`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
A5gyKW/TE1BLZ24bmmsl41T2LXoh7m0h2xf4g9IYfE9h4rw8O79vQ+NUQepjluO6
7TA5NK02GRMS5mZWcZ6DzUNIkSjIHWfIORUxIo3Buw5Hbhpzew1pappKidf1jqjr
v2GUSIxH0/JD8hdJmyZ3nP/9zzryLl2jjFMZwHZkgJGHJF1cNfok33E3AP9GPQcv
9aKB3Xz99aqvMMMPljpEy3FzNzsdURpAyY+irBA2FfDh5s8xaP4GzFjMC1PU748M
j9/CCUFHKlhnZR/hJrCWwAnOtLN9nLm1e1cv59pf9Lfzc5pbJqDgBgYSExyAyCAm
PIvZ0ehE5Wbh7EiXZuIMZQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 576 )
`pragma protect data_block
Ny4pB5aybwc5/AhoNzITBjb4cRRn4MqPrsDan+GClV2g+6bahwNqiVEHrNx1/fHc
BQGPjyY6RSpEkH6d520ESVMI4U/jaCrYKOHfS3yktEwOsj+mM17edE+zJdaf/zKD
yCrRy00C8gpBMOaWUDFcSeUVMTx4KDt3XyD6num4qX87nESEIyIbEtkN9vETeXXn
n3heeREFCusl9piKtdsDZ/8kRkgG9IXIHb7Lv+3k9bD6kVDcWl/Qg1qoerKVLpoe
9ofJ+UW6nC8BhZCB2hVDBlNdPddCbrT2E3aVpA3bptL7kLDBOI20BJqdobF9qUgo
9si+8mntjb0UMQa8jILVYc1kAh3CZCI6H4TM5a08n7LugavnoIIswDxjrYvf4J97
MokaG6QGG4XZrtVf0We6JrefLrMdIxVYyezSGsifEkguxU2YoFmfYgKLDTlCrs5d
nxVX2KVdk+YFPVdxJkZ1uynm8K9RvbHeO9f0XkBDT9/5ZbTfzZpEsF78SftiJq4l
bxHGWXg2YNrZgs2vmcEXBPLqzDc6osgWj55z6DrmCq/eflJT9RCufO0dRM3WAmri
jziEM3zuLDZx7eUxSR8p3YNYx68s2Xl4bmwI1pkZry+eZx5OscQyMO7uBLCMtOx2
oY3ioF3m3ZgsLMQEYrAzgwGjjattF3lMGciwAydA1pnMekiD0OKcqXO9Cf4Nwazg
7WCSG/ElxrwuiIPKgcf3sZygpANr2yZb7HoVI2DsLUK7ft3zamEHfed9QJORkZt8
`pragma protect end_protected
