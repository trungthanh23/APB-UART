`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fZtevKrr7LSpVpro/vruJ8OCqXXNtRteJv/+g60qicljhMkrzZ9oXGtxb2ORDvVZ
VAJxSzDVAacPfsUwLCpMfOyMcbhQT/wEXVn8NF8xIDuNFLmkKIB1Ahftypa4BT2U
eSKmeU1ikCZ69olRcSHC1PTcQFzD74f1nIedX0PlBbdWlo3VEs+kGdnErkyzOfDH
pKe4irvyicWx4RO8CgQokxCI71LuYKS0yKGElIc/5kxAm/aFwwZ1fpMM7LZUIIik
KwKl/yyg9Ec1INM/HXjytd2vf83L9kYYckh1ve8A7o6w83b8n6e+WknsSS7G/nOF
wcmDBLqJhNEqXg3LQncJIg==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3904 )
`pragma protect data_block
WhWVI+kPw7A/4ii6LCUD6ob/CxC9RkcN8P6pyEdZ3WZ4BLJQDcp8NXPSc/KdQciw
9AUyyWuaNCwVphFFH9MthQgvE0AEilyJq63YYVIQTk9OBi5Y5OrU87T32GF8DW3R
2Z7o/h6RiAura/CmAbti7HspEcrIooxdYhrrGNMwJ6A3fG7rTmTH0IRzgiOQKqjj
9u34WT/nvyA/CNnCqYStSzfcJwc9KTY3St93Xhc7ePfabQjxESim6wPyYTMtZmVO
hgGDw4dXR8H0aVW9x89YgPKjrNSYN27x3v5bMg9XLJ/aUmakNoZBqCAijvh3STjs
pEm4hVedYyO+y9FAuQn0rlOna2qBkIOAVvsB0gg6qkiB0ooQjBYyOE5d0ZLI0oSs
2ZgFAfE+1pD86ScnoDlQ0MrFFqvgr8rOZ5v+gIjJjn31Lh/r96U8OD6EG9BO3p3q
T1HIfz6h9Y8lljh12zJx/rllZroD9/YmftzDw+CsWiQVCe+Fx/qp9nNFrDmp9HhG
ko/ADovzy16o2Hk0Aiwaw9hKB32ETJXu60J3rJlF1o/kv9hTUaYV9eA2VDVpQEvL
HxK8SqdKEwDXMT96Ed7kj+VVsH1uWrfHYdH9NL2XqqtpwUX7GRfM5RDEW1ubB1k7
mF/Dn+Gx9J6PupgOwPAQ5DDsH66eGCHmHFaquJQqrZFRex7IDSmly+JQ30Gv6xOe
zcVriseo+3YS1SpnHzhXeYmdstaQiZrNE29kX/UhKfQM2j4VO3tOjT1Q8GSy/x0r
MDHRBNzZY3w/ASmNBbg467ZdSbUZiDUzYnUvJHc04/QdA4+D8dtIlxXVMua0UIjJ
GcvNj8VGW3Rgb0Pnfpd4kK6opIEd7Z/PR6j7PYfpGS4Qs2kQoNp8wHBdy4MU/pbK
7O+K73b4fLPM64ccDRpRFECGUFcEs+bepEtUPt7uxAkWzyWHXK7FrVG3X+jf0Dl9
qg/RHuOdU2vR+gXG2ALErIqdsplykg49Re8KwzB4w34g7rHKatvzKzLoRwO6/ilI
cqclGDlom1thYJoIYbyH7z56CjiIMOCLmvW6lX0s3Z/FEzJAfNzkm/n1hBCndAuM
ETTrR8MRMybiRIbQNM31QOuxFm8iFC54Pvqri3/038gx/cM3JCk7vwvg9mSCXsAh
nBngkSHrpNpZQB5fAnadQdpUODxYwY4yvatIf24E/qptZX/TUtpQnNS3tVS3Zg0B
tiMIHZ1H1BP4Gq7ol4BRdrGFLUbwVkVOb7f44jS2FTJhfwQbwoV5KlYKn1AVUhxe
z1n1XxrEh7VaBJRGTSFwLSuz5J22LOuzJa4t6+T7ugjFsrV+wSmdZ/njYv0cmzOK
SSfcPoccAeZRzUsBzBtijY5eRHuCVIljecHtKTf3Gb5VTet92npCmxEaJIx0iO6E
CLPb6Om5026vAzZKm2+qwHPwGttQJf4eRXUnYglPgO7QHW19MFce76Nc+hkLTGRe
xbxZylG/FcWY5EMeUlTFZQMDZpiZmID6JjTCLkWK+twZaR7/9sZaeaxyhyxS5vTl
V4lcNBbt5BWUJ+lbyR3mzlDzgy4am8x8Jt/A3HWLfcxtqZjM88RVpUPlUvJNUBOR
Gip+XDpQs9pssz/UpBaS1D/H1Dsau71CfypOWV+Ca2uqpCqEJyCPX/FXB/HcyCNZ
WPVDlHCwPQTyH6UeQ+F2SBOOt0clb3pWW90G9Zj8DyS1QVXxcfEcJ6bPdlk00NUr
8Psfm7wHjTcII5BJowV+DF3Wwdf6J7Ebp2TDAnhhXGW/fZJjB4rgGoxOKIBhSaH3
PmJjhgsJNBQC6br7Ij+ihAnIJ4b+XFnSscD0LL6x19YLYcjyxasnm3xQiocDtomA
GsIw/1QyOsz/0OMp2nHswoKEaO0xwsIfjXXVqbZYlEqWk05Io3TMV8r/IYQbCia+
Vd5Knk/EnPv8YZrLxS22r98l9Kw/vp+8WkqqnZdHjxp6gTms1kVHtZblBkUIPLqy
0HtOzw4Pugcaf/GC5qZyhtAx2j9VU4Io4EIZ43b481hdwr+tL/c9pAl1LE4CMQr6
wQbdL7Q1v0DCU8nNAZZUjZiNQT/5rrE9RSQE+4jb21lRO2AloGSjmcSrSRsJrHzR
XUJ4evzf1r1nF02LYTbPavovcV7KUK9ZXB36HJsGydBbkCK0wvV5tTiPqfT1h03K
ylpr1mEmlk8BOKH+WLG25zzkkjXqdt8hZ4t8kaysqr7juoVJuexgbYUSQNQpMGYV
KcbgHGYwgbDsUfgJl9hFMjG7zqBVQMLGMfFniMF27pL1zLe83T8MyzSfpwJ5gKAG
wMkvfZWl+DPSHAS9PU7O+RD5Pz+lYzdnsoucEXEMPc4rplNBV1YVAIiCAnq5sPgQ
YudlqIYurh/f6VA6LAJ+BTjt+FoWydLSDk/Zkz39ddFMENiL4YA3ZT4VzL1WYLOh
9CqFPim/FcMdYRF1qKACxOZ5rMuWs96fParamSnsYIHjkbiiA3JlV0eLwDpjnJlr
LfuCpkP6alfUVmYy8uG0LTWWEBvpRFbb7TSatc3cTH6aXQDyjkokTq2ehROH4GGp
3jWsAJTLOue1kBx9w8D/kLJOixb/k0t4vMA0sj5SRBtMtgX1yEJRUgqUkEB7Ts0e
SZ3xOGhaIyAnnEa0j4GsMUBcIYuLpKZzNFXC2FnRyw3GksEV4w7ccsW9+RSRFebM
NGWtc1LKkwoPXpdY785irvf9XAUOwhI89l6QiB+IvQ20Kx/Tnmjkbzd/6/aPzO4O
bS9W0cwx6n0TpBmSVCpW5uMI3UgaEt12SfcUw5jfRboLfiFj9Y/MocKs8CWFQIco
OsKF7zLNPsSDHo15N0D4l1lnKjqauDJzV6/wWQDO+IDlHPTzTJ8q4cfSlTdVv/yR
qSfOuhko0ql3U+3FFNxjIu63IWJlUgaKU1XRCZYJ3hZ6bVlViYkuZt0k9j0hnYzo
+iOLAxIEA9xVpPyAmlMrcYEzgYu7AYV5zlHF8/9TecXN4u++yMzqKnAoov7CMZqj
Xskp0Oli4x07mBcQ56oPHIHRLyuzUBP1WsWriMCIU1zo7lRKLkudVQ4j+jfWOGK7
ncJByNsCP0O4JOuz/5mCCCB8Cre1P1YFIIJmq+JUnPtnAoRg5LwG7DK5eyvVj5Tt
c1ktdSRSIgejoQt2UVvTDLZgkV9JQiLx1yw7qzByLtDN8KGp3tnnGowjNQUZWZ92
XyrXUTB14rw6ub3ccOItBXNXZJD/cZmvTQuKBgzaoU+b5H/NPmLIwMoxZy3jDbzu
RpQAyGf4BkOg75Mj3OQMxs6gSI3JCk8n4Fpg/uUfKk8Hx4ReEY3rKSMZ6zUSGuul
oBcYT7bDEr3qN2LzpRY8xeaVzDkegkk9rw1u+wmj2UEH0bcG8ULgPWFKFThnlpbP
NrLmlCFUST+gS8u6aLE1bily1DtBPmZJO8h9w4MNpc4l0hB2OMm3q4VbXw74kJHz
TULqZlIvssDUYiGKReHUA9MtzundOo+WWoP0UtaXkCpB9x51PhMNngUdzFWFSf7c
pNU9upAMpqp5l8g4I3or5Gm3Tj9imbRIbqn7v97qcXt6cCHiiL1bph2blMZwtIJF
a3rPKVEvACHhF07M0NUevyHXqjMSSJobn9QltAQ4f63EAJPGBriSb2RLfc+gat6L
YioNbyQ+qD1ykJRMGs2YrOFYvnExbAYkOTm72rxeVXxDgxhiRPTkTG6Tcs4rN6Mg
1+nFd3Q5DpS7rH+C9yfUrxUhMeLUVTLx0De+Eq3S5dyDXK/u7oR9FkZcOZi4fAaO
8stsAD3oDu2OSamD5vmXWLUotzU2Shz3qdd/kN2nQ9qFTHqrv/Bhg1BylgiVHVSF
UKJJq3YBoEegtIBhSkgYJ+E4wNy2n5wSvNV25QTzxpEul9Pj8dycB2Uf2eA7OYD4
Sc8go7jiqwHG2WsOTpJzeaq2KktKmM1OKguCzjQX8hL0NnuRUOECq+IDee+bUAow
7oH7HvlQ/K+46cbzrLV6meV6b6500UmNFht0CyXhTl+URnVvsi9S2dXWF27B0ral
+1uZIr/oW3d2sxmGgFANy/MGQBXuHDA2pTZfhD29LS9ItreIpBXFm9yGa2N6L40W
MBp9djxub7va/UICz0qdCcTzIBHsyL7e8H+g2AiOj8VZV+KanNam5nGzFfaDh8Xy
FdxRwLqrwoeEdYwDTINwHf+6jorNDkPunHeOctTI3TZsVVrVOSoAiX/qPt9G9tnF
QgaO/zFfmrgsQFvgS9sMWRa31munEaPE40jDmhHrv8jgMtqhRPNw+Gzw8JKL7P5t
QUycU8y+AA99HwnzlXgyCpoH4HI3QGsHeBS3XsT0vcZyI3XRbmw71dqvqhfeVnul
ztp5NT6c54VQN4Hc+8qyavbHr7FKBM1XJQy8GY44LQWipF6118zpW65u4ezem2zz
gHKIxc6/f1vm47DXJaE0wHNSbl4x0ggYa14+8CKr9/cyd7ijrQ5lEgytymEB+ygQ
CX3Wf2wTHWb8AaMkY9OPYqAWpQ7JsOtRC6V/sSVQX6KEFRExeThVyT9bCBCbHIz5
asnMOFLIx3Z20qX7dpr5MEuUlVT/raCtaCxXByCpGSLqOI1lid8OWTn95oq6BPoV
IDsXw7ZaG0rXqcG49FoPIVgJHvu5iwGxuWinYJ/xHD0Nz28Fq+GTqOvttzy+DMh+
WMysXREQu9FnHf3EHQeTALo+DLV5G4d8a8kn+ePKk/8TSY6lsFhJza9pYZGQkFyH
oku5m2BWakcCFxudxjf94OBKSkG7uf85u1kovnOdLPHBngUS6kUX2dZhhZOYs37Q
Q1O8L8fKpMfooTVX9cRS+Ky/Cs7oEqnlmx2xUguGaWdDzElErqvHwPaXGaTHux6I
1CPInTooMmwEh6jfjgT9vs1rb8I2DlOJqLZEMRj/Ww6293tZUPC0qAoAXcK/X4mf
sl9mAYZvc/IYkgjPHO6lgu/YN2RRZLj30sGJNylTvOtZFitnEyZFTMjpvN4Ymz2Q
I9Sz9qPB9xRro9FA93Cm01nDL6kzBpubRaGaLOE22DxrvFdMwqbfQXliMWKAuZWU
pVVREtgDSk7sh+Mf7DE5BtvwqaJRnqoydJDtBU4lUkwy6MXvT6FL6jQKCLt2MXuE
/lzxk8aRhQfjZUcqHClGiIspfxbU2aarwUFXqBLqaGxOF72wNWACZIM61w9SZoZG
hBuRKv3iXg5953UGV4CMnA==
`pragma protect end_protected
