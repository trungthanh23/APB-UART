`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Xo9bSND58i8xrfyJEcSfF0vZq124tDHV9umpIm+pgpN9wFz1XVp9RPopf1+Debep
95NCbAfOO0vKRtLwpkDx4q2O9ouN1MPCPJH9zCbitw05HdvjsUy6XF71lRBYpHua
6YxGWzZuJtyBM/NU/4CYhixPiy30ueipZBdx6CK06ZCEZOqSfmlSDwUIMJZ8N7UN
CqNptPIHamTQr6fUludPLAMpm0JnyYqKG9uIJiAmV3LH3c8cG86n4b10mSnXweg0
cUx9rv+oFv7ccK2gv++3w9MclLUL/yw68ZmGG2VzpWdKEDhB1xTCARqsWHujzT7o
398i92I/pBPgnIhPXZlNvQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10192 )
`pragma protect data_block
EkQH2/646L9xtAV/ES5U1rtEbCpJk2YCBeWctwk2iZSN8glLtiHXxoI10bjZe8nd
4jdMvrtOi3bpwqKCN4pmyFBk+aJb3oloNqJovhrrSxeB9bv+yEF0vRYAYiOMLVqb
3Qh6e5WrCl7jPoM8ocmIVThEb6AHpWux29LpO6Yp5DJXUKRmV/qsHgLGjCr7rRt1
gr3HADVbMKWAQonln11JLH4WQLvhAp8C8KthRzYKurVT6EskHsH/hX/z4Ow95CWj
Xm/xWOXHNzoRdUNb9RAnqAYKI4O22LXLZ4z1p+TZNkLI0qcjrhoTsHNlMnYjzlrX
hgRm3BCPiTx1yO6uCk4b5s+EU0QzYHt6UZkuWqgAkBLWLlQn+VvILzdZ+255jmoV
Vxl8Lwr3qEpnLqP10AGSgRTo/6LFCkaEJXG/9ccWdQxsWCBlhBdwoKeVLYijMcRj
HeOlYnbNJUiW835jZJONBv3jOyn5hI0fZX+z9+yBOtJueAOQFtOAnxPiEew6CDkE
oS/JuTlC05LlovcrEAGW0s7WTKYbDB0Oumun/NPDpH06SG8cJlYfd52LRWv/gQwS
/0eerV/caiy6QD8NZKnInhV+kjUyNtXGRqFNhrD6AZHMKTXGIbwf3aP6ZtVZcbGg
ImIqjRAW1ZXRKqrw9+3tDUeahInmr6Dc9Drkfv/2K8nw+Esafp1aiOUTdbzUgRsj
Xxy32ppgNRywhhkGLwTqF8PSqsQyrlRZXF4ZOUKDjA1SXDoq9LRApfkc4gg1899M
4hMJRmhPIXdZZMQwDnabSb+T8rHM9T1/wODNDMN0SQZFS+gCSDISPI0I9TIY7awU
UoX0wEgrBrqIA0Hdy3i8n0b23r6Ae1x9ETiBEFvJUq6Jp3yFrXfR0E/b3hknMGES
DY6Vd4d3yv8cdkUSbLYlbJ0PL6ysVRsKWx7ERiAVnQXwtHCwZMpyxSRDRCd1h4QK
7gOwqHk92VfKDn3SBryNV9Jl8Ak3TG1KKYiZa6e1TzKiwmhb+zZ0moMNqnBl93II
UuiPxTtAbI97eNHvJnLICruRhOyUv040Ir9NGKiMZjXtonuX20NE8YLmTuTPJ/hJ
VHso66kRildziKojyv0vd1zzTpWQ1gXDdGMrHvKOiAW4YRmS3rS44yXS4Xhcxk6n
3ZrYADnjL7IyuKQWY/Ki4iKpL2qnzgpijtWzLTws4TkApDIS221PkyMb10tC7mgP
UecZ+9CoZeoOH9H7xmp4jatKpuJo88r/QjSYRGp27kUAwPfZXrcdFEFLJ8NunEDQ
/m7X0L3mrZNyTnruPQg4DrM3X7ryyptPvAEu+SqdG1Fe8DCaO7trmSo9ehXE3Gjf
ryxvbrVnQxbbChZBFX57UPv1gscj4It/+rRbF5CaOJ7Nph8f5EjpTCqJyCWIJTAT
ue+tLDb04mQ4w28dG4Xp6ZuPa1hFToM/0xTq02z0iw7HlZdGzrrrJjAbS5KPHp0E
QXr1EmcXyxRMsE6ANeqpnJLn5zu1VCAeNVpTAmCqHXjixKWXXOXNDT95fTAADC9u
7vc6mVgQH5rKMOiGrJ3SIx1O3A4dh+Al+g2o6OaCI2IQlbBeWcpU4T5aYPKUQtaw
r6xDFQV24Bh7s8OciA5fgR7RMnPL7wfICbWw9exWgbT4OeuOp5QbaR3LJfp7c/1O
Ef5dlmzZoun8CWx/T58RMuoyHDiyZpelIxV9frn5QZH/auaDWLaX9F+oL32At1Hc
ppjfU/zbNRHmiPkvkvlBb7G2gbofJcqhSY1TL4xwGJPzdFi36vBry1Ms41jC/d4N
I2omByqWpN6XDRMoo+TUl+y/o7ZqrWpZlywIc9gGMslOYR1PAZYz2K02Nb3UNvm0
Twfil5YUBNAQxzG4NkGFWC3az/mg5RdDD7vrvpga1h34Awhkit/zxI1ze4S245dD
2QTQdrtYJLBBaEqiMQzcJV5JPJTydjop64xYOyqrDXCk5kx2BklrNRPfbe792Paz
8HhEM6fMX7QOj45se1GQ+bce2yHC0YrPeYoXcGqj5hewQ3GHXJSbl6sEaEJYIxQ5
uafayCZGhHzDrAmXkdzskjh152pTFM01TFo1d6cc3Au4u8sAgB/j6ey+lVuG4Qcz
5pMdbpVSY3Gkg4NqgumqbNe6VAlMSeHGW9uKzjeomtGlwsHu0VGFL2NdIvL0ymhW
tULcjQ6Uiuvtbp0CQKmArnIGWleJgZBjUek2ODIWw7GPzxU//txrAL/+D3fS8NlD
Z1PhY4ltihm9z2XAFdoHDShsiHYLZcwHl/ZZ7ORGOBN/HCkC7cx3I1eqnaBlaSOf
SvlF1nZgHSekpKaQ2AvKmVRpoO6xuKwzC4thA4q4ICdwRIFrx3m2taUgOq4puBat
zWZrdXF5ENRuEPz/zt4t3ctIlfwI5q1B/8AYZFFxBuJQE+fjBBpLH/xij4vEh+07
PLqfZkp/d2nBkQ9wd0o7YKzG97Mgs9GLzb0SRCBHjxmIJ1OW6uJRhzlW7BhN0FJa
f5jn2a1zsjCKxJpV2bRz/VyOL6nRMd5D+zcyR73ZcWvpx9kw7mG+GaAApNk3g1d/
tJ+LITdr5RdFtptQVLEXHeDxoHgokoHf/hkQtYcVkbVhkf9QPWFQEbWWHCnOPnKn
0Eyn6nJDx5CBWvRoBdTbU0UM8DaC+qEDzA7OCHs8pepefzF9UzrWlA+xNmFhNs60
KAYhsgNukH9UTZIBuj8yUmezL8sy6tNi8N4NW4U/kr1PxZVgdkqU37TuRf56JAEJ
/8Y1C/dxSjWtaBHWf9oPetEA8bK2exAG/fQ0VAFonwUSaaGfwoZkXBAemXv3Y7mO
cIJSwGGeZmUR6d35Xyvg/ISnqFlOmV2+tZNYUdgO3myjpomalINqoebf3JyX1/5b
yHcI0ddHUPc91eAVpYb2cWCrFKvgOGnKHec2/tmEVvXAnLNeAANTLsRU/IbY0q0L
hlFqexBl9mGjf9sjGn18atctrIw2S45v4LpEqFYhu52D2vKAnsDLG4g+qoa43Lvv
bfX6oo56HLqc1z8xA8YXdCkRES88yKHdgSJzY4nqGnSpZITSgme/L5/lpcS/zokj
gJELRxaku2HggGjKzYEuHwAiWGdafFcDCr+WU9ONX9fBYwJ3y/EhBAoqhN2BIKhF
nHz/qyC5eVJX3pT1/UqvYGloz64Ua9V2GFMUyZVVf1LQJI1oQPKWmKrkXRPdq43g
dxLSbpdqPCDfQBisl+j2yJy3Bkq9sq3+GO0NA/4vjM4mI8zc9myw20gMMOUO9D4H
3Nl+RCASCcNk2olo4IzJwx+m0MC/nz9i5t3cZJzKfItY2aDl9EBe6neXouaPORTQ
rTEsXD7G6tQ5vlWEXMz43mBqiqv37NT0z9Pt1FcvcV8kducdpHvwA+khMntUZrnd
IsgdyWBevpetzTLO7YJi6jxr4JoJDcyZQGG8RcsEDCztP249H5lccYbYiGM+K/G5
J2DBezLc9X7TebdMITs+T4GcL/fMbFvZEdBgNFisyTaF+TsqOxYxjoXXUd4qHQmf
+1Pyorr3Ni3tOHiZ1vGUSp4Mww+oOG8PswLYke5J3du3WAVUCpz6yo8mbSc7BUjG
xxtPyrmF/C9jGaj74Go1jSPlL3syxnkBbtahuylCN/ol1AmLJrXfMuX/CpHcYDDT
x3Pfqr1T27THRVrWjm50FXpdcWMBJvug/ujc7jtQ4U298hy57BaS/sN4o0+CR1hc
jdmQCa5kvTCnEUKtXNmL4z/8Ylv0FTh63iXFTyv5JbD562ADZuyBUcbmzQQpJ6M+
dhPc/mnCbt2agQMvrQ4EofOvs+SIyVz0eXLEfd7M8IUWZ/6FVcTwml0AkDKytyBP
oqJ0+o8+MFROppuPhLRzqyaK/xTyglyibGSLb6FhKZIaUgPipjmjHV4jr80WbVxY
f7zCq0E54W6YTq97fqA7PfEjejRD5KGLzTDPNSOwsGrrThRWx3gswkBdKNnlVfvY
b9OomXKBD0OlhQjiKIMgT61QwD0pL0dCRYXB28eTfmtJnNfyQT7bRTGAGBwNHta5
fQLCsL8fnC2NWGFrLvxE+oa1tkMhiL9HdEb0cdmqVRPj+CDpcCJggK9zC0UDWEYx
HP7Coky6x/lXOKPMfxlTLO1jO/lyejQ3YiHiOzyvkp70sl/7oy3wrropHcXNCCzw
QasGisYlU2HdpOaIrOyucUpnpwazYfV2FSRj7BWH8obs7pWbQ/N9wI4kbOYtYwXi
J8W93/M0HA5o6P/JKlE0Y0fKw5xvCQ4FNraJ58WUNfgULj3zg0Vt4qVTmG5YIhWW
PNPJ28CQZTK3B6COlDekHO/pa3Y2TmZ7baH0y0kNTfveAAg+ANOb145M38p4X9QJ
W8Ih88X24YMQtly2G+anjnrbMInW5pufPkzAe/ueHFE4LpyAMpSXl2P2m1Etqj/l
oHQEyiAxBNUD5ZUvDAe30IUq3/ui2Xzn89khNKf5JVEAICGvLlv4EG943EUHe9f5
zXmGfDCLZeDi2eWmztk6DSoDnUDdUjIuLHCC57kn7h7JuLW6O/2HmKImd7UJ5HJD
UwkyY8b7H1kGwDoB77iY963WYQ7MODzdvVMqSo6FNONVrWJLQ8BE1z83NWM51lAq
lRNe9dL4/sEGN5cHHlIcvqKWWHAizhpKTEIREGvHrYY4K0Icpj9s8ve9Vlvh2f+1
YwDJYxs5fw8aEhOEKhC6z+4oexOOGwz4nv5I60PqyV7z/dE56wfagyw1fmuqmnpK
LEk5dNKagA+FVIhIUVJrbjryDllNzXRvrrjook16Fpg47vs0c3Ie5f+g+cYBtdMY
rxKIqMSTL3JiLIeH8H+rYhuKE2k0xc/1zNfgSgtVkqY3Pf6qJ6dAs2wwSFKzrJU3
31di90DNC3+1ph9adro3EYT9sEuZstxK7zQA0pYeTFmJbNWPjg/ZRr7Ba2u0n9j6
rfE+2WgytqKzH2zg+XHJn6zGCxb3Zx8g5n8bfi/8NRnWD9ibSlyoA5zQsWPefQ05
wdTtlq/GI9Clt4nklFikVoPoEoggmiWPugWjjfKc2MZdHfKhWrmpQrOdpImJ6eOg
/S8jjfBhH+efVLN+YQRo9zgiKFJYmIcTKomT1UHsZxV+f4BA4i8BvRK/QPg//d3H
R7/Ayg5qEbabmVT5UY+qyHqPYOtVC38dvkt21wGkoPQ25192Ot4k/MJP0tmWWBzr
3NzqQsrYX/gV3PmxfhllzxXT2tU+ysIn24KlwfVdIhrTyEiPitgQPboZXdnmteEw
4HGBdqMG3xaYjJIy0lo4fG6qizXig2IVp4VjvJLtf69icb3p3bM5gM+BMAyQ1adv
RjB34mpfoU+3MycJT/+C2XgT6w8MZALQwsz2JXvVSJxYAwr31i1hoPucPBmKgzwM
KDPhezlOTpGIApVfaidEtmDFRLJLy+WZsVHeX4EwBlSNDjV/23mJRV6RA46O8KE3
ZTjvRTH+VZ43pZWmmZ4i20cWh/D/YaYJSvazNZPh0u31X2Ie1NObY7D2jbAjeCgk
M8uAA0Ujq5A6nrzQ7WlAvdpg2lzihS6XRgr54aRtP00kU+bbeZrnhvgM4cWBQMiJ
prBhnEsD0+KoSGE9kjcYc6DcKVGs8Tqh7mieb2XXmPHf2n5JvRX9sLgemvBbS7yF
JhITmdT9iTSPuzCLFNFLCwxONFK8e9hNgt6DfTadqwL5K3QQK6/nC/phrYVwJ0LX
c75ADA2+O7QKpBqYfYOOdxl15O/h0LSqYZWxcWx3xxpDPhruet4KhkffCkbE6btj
knj/70kTavBovDpZw12WV6jVfOHz1bcYCzgj80UE06IVLM18s9BFfgety/PN/nFz
71N3IOAOMH+Q8xuCqRXR8EHzaPp0Kk3na68XMADzIAG5ANtCL0XX1p5KqDBs358a
s4Fau3gAeYHObBH4rYStQd9RauGp2B/6JGjdvQsc2IfYEdIGYq1a5XwPAKm05fGK
8z5RiyHg31eSSMMwpagFXO68p0/cSbELLNYUxptktVNMM9lA+GMIJNs8YAV55qI6
VQFStgYc/SMkVWE9IWAtmRuqwP5bFAwoh1k9Vx4jSqzRlYeUgG4/Nwsy3VPp+Ytk
F43POu8p2M0El7+NDRMRv0rRDPlSoPIyVJ6mmPUe6szKS4/+tNMDh8uYU4NbKeDs
99Rr6Vv8BA78WXjRbj1zaXhTWnWVCEajI5ulclN7zh0o/0L9ONM0XrtSHlVeHIfU
rsjh2qiAFLSE0ms8jnb3yr6V7S21clPNoD3UlVrQhcT3cdbsHePMwmR2qH+RiUNS
x8OFQKmpTKElpQk2rq/mlD0HNQFjnVUtnewZDDjDu1Y5xtSGKir3emVf5PUX6cCs
mpVg4AaC8L00ybfou8iV+fZRbZc5RZAaGhxmh6x9HTSQC0QRQdWk9Z8twaElsNbA
YQQrF8POdfRm+56Ho1ZtgTMOSuhse875OxXGsBVq5PW++WqF+9H+O3zCNI15ARDx
joFgFtZRJLt9Jdc+mUA1J12TXmR5edpRcig+3vccYG8miSXtbrUtzgRj9rcPiOFU
Oxnt5q5mugtcOJLgZCYiBrUUjHJcPtfMRGt/LVcN7FQlvPSIIRpLIwsF6M0UaXfl
Zk467GlEIXupT/1JU86HcDw13RKN0LO+fMBDyC+E9XnbrXiPclJfqvOdYfL4d/vp
gpq1Wz+KoeDI9qjc5IlbdqBsAHRQL2nRYs8Irkw3lZyHjTu8b2kNpH8ifQS7CdJx
mqkkPyMtMebsQGmbaN0cgTnuvqMjx6Xt34ukEhbcbWCPvXfnBd9SEpINZsNzvMGc
t1SWJ/u+HHovnXO2DK64dIoI7ckb8Lzq8XlEOzZRFjzW5HqXXPGfZrXHPVUw4Jr/
5V88J82c/1+qy/iAY92K4OczAHP7A+khOTkSw5t8AYIEODHNjE1PpFbNz956nGmR
ROrAYBdofA71iqHEeVeHNoyXq0Tg0FnhEFWfLmTlnhIAFdGShDX4WgmEegtamr54
rc7hZVKFiF7sQnTEd8WTGnKxj6Z45ewJSl0V8fxxc+bm6yE/2CVQS7A7aIhQNOqg
hXCjVoBx7qC7L13puXWfTOdCsjEuVoBneHDaEMFRpGaA7iO4GazTMAkftutMLqVh
8yMgrWHteH4VeW30YbqPoVxWrFna2kIXSxQ3goibB4qeEducc3JCxgINAMKd/yXm
3lf4daWK5wVtxx7ZBqq4EpYjHF+ugviJseny4ijQY1AfemHz+U/bncHkwByPcDxC
YGcTnaG6F2fZaLbrfeNdU5MOnx+te+0eHXzDPHgPfAkyHM6OGwAwKD1ykFjdlh7e
A4l6qUaWW0TaJpsZQj+bfG8xFXZrSUMJr1riMeaJZvKhZTeSKCAEoQ4ID7GzAWV/
sC8vM6jUp3iRrbKvdOgYemplXFgVIldcj3Wxqxxd3vTOs0Z0tbmCOv3xL6490DMV
OBiHgomF5aZIlxiwuPfxDCSjF81vCU5W6aBhtuAJpZgF3FgIwGGt5cznVlB40HET
zWgT26jrvt8QCb2BBMQXLGE4nfXaxjxJC2rwf95H+e28TTN933K+aQW49gX8dU6W
EHo0AxLNi9Q3YBc/rHMPtBGae4sWJFUoWpx/2aYIW7TAjuJIlV47hsFaNNzZmyoQ
W+aONhvl7IbB0idUP8ajznVaGmI/mmLoYJ1lIrk26puNYOTjKuXwhT4lcORfv43P
kvktl9MRfW1dfcxcel6/HYGi8wx/sIguoY40vN4oFXHd2cEKjqw5nM3ZEqX37Upa
yB/EbBemc0uD3mfpLLDqfvjaR6l8OUfxQekfXIxf1odMudUijbq/PbCvljFVfzwb
Z2EieJcbfjr/ktcP71sZCxHNrhcLUJ/YgkQhjRvDWSdX+juwXUwTWHQLZ9g9nysw
u2AIDBMnCkCMLDh5hSlWi30nq9hNjRv3VGTF0NGOoGgo4tDgYj7+m9s23hhhPInY
GnYyNptfmB4Gai5tVZpT5mDXd2asiJfq3dU1+24V5n4Vim7jYFKb7okJF3lvkB+n
V+OjE7gaydM6Zn+JwRk3SidMSiXWqwKQEb45yrjXorWgm0+8KWekFhSsbJLQuPfI
oc1+aQ/AInHoe/5FIccjg2kufvJCH+jNXzsl0b7k84if6GLmKz9W2fd4yJjnBGxv
HPQFmp3P52DqOFBatKjbmOWlQhejqM0oAJ+HQmFsDUNP53HTT4GwbMzUS8996u6k
n2gpRNjb7qGGeG79KI+3kDmgTBqBbojDVOiMO+QR1zz35wSoji8+/GKPhEQ0NM0g
Ww4e814B0UMLwRV/Vfu29Qxs0mhE8RHzfHXnBWqFnoNOTBcCxLr0UQncg72QvnpH
L9IYGFsZmprJYJpQzjI9sWVwtTjcZIJW/OIU9+kP+gBAhtPzAmcii0VFk4s21x4g
0EFnUU0V+/q1CJjjVW6/mgJZocwvOECX4qkxQ8UIcpwBZEiqo4EUJ9aI2cgX/6au
YrWidjiZkVfgXJ6o8SFoDnfxfUeX5RK3QwxTAU6Rh0Xa25wQwNmCCVDczpnIuL2e
YpcgzukNVa1ZydNLYK/2nitzDxqyouxKwwOYcFFkpIC8uqRbYDj2Vf7QLgUwdfLx
1pE9fQ7/3IIdjOeU0uIwMLdvAoN8d6DyH0QuzmL0TAWSXqDap2SAfgBLxnuiAMvr
GFSbtlWV7wk0+0biwmJRoa0wXMNfJIIWhgHmCfjEUou4JprOrJeyy3KdOlRzsEMn
vC2r7HUR42Q0/R7p5fjIOBPnaSyF7CIOUuFyt0oVooSV1GzRiW/CGS5kRzMc+wpu
kRGiSIUkpX7Q1vZWgKkR6ypufjIY0SvuSw3RkSpfffoTJGt3lEmKPBqKw5l8NriF
cAg6sOLgAnUsONLOlmamsihi8VkIRXP45PjTPceQxoftUtjzPAkhsHeREwqA+N3I
TXZm751KcqITuKdB1NBxJ5AZNZb58a8hmh4yILoogI/wmoXup6uz/Oxj2eYOKV4b
FkGsO+BcSYZ8kYiMX3FOkX5evFSH7JFb/4tglxwKzlm+OdWN0QgV44ZoXbyEAt49
f8vIwhWWZAOV48VZVqgWs4zIMiMwlDZymW4FxkaM2/zFjd3bJ/b7BA7tJlYY1F/N
X3rNtv/dV5hZ0eNTNAPgMKSwYiBxs74VGZ9Ri5kGxYOpyNUqYRyUjR2d+ObX4WH4
v8rfzd39lrQyQHIGgAn9AwBzvyVoStue671xeL5bOre+ILEYbGATb87Wo4zTm9xh
Ban19PfvwwhwLtbXKT1h9X0lqSNhlPy6N1Fahrte9yATRSOxZr7FVl2HX85G6ecG
+pn52lpJbhULxuUnZ9CeLMpAJladBqzPeO4u51dxSu1Bi7DFuyDxQsyelkgsp1ln
D3ro6/hUu9Cbln1UuUqRF2RQDkuNFS0YIz/f9lFYm9j9+oRAT87p5G304l56r6Lz
RILCic9gM2Bi21ivQBxYGK3KFbw6ajntmhVCqBZRNTATpFuAe6JrO2wkxVXkiarJ
2R6iELUTA/AlS8Uf+s9w4CuR1wqPuMy/QcGFmYZs7KZaT4ys2Ox0gALIgGj+3F8R
+2gJZUcv1xLFcVZNV5FgJc+DGIuhqgZESvyWKhCaMt/d6yIvCGzmt0aD9ZPo1h89
VjkOPK9gEtaqNS+eKcb3vpeTSvjyRPlfpYXuVuno8lo/Gvtvz7CtVeyhWXpMEwrK
tq+GiP401rcpDHZUc26jBmiqUdxNFTE0zngT/Ft/qwByxY5cK6VE7g+TpSeLDUuu
tuk/foEM6BHlEjBstdkNzggq0EYlMM95dslT8812yNLaBsJ85ScScPFYRocaftDC
5ZuK5bUY9qntq4xS0aUmdYXaNbn/ra0W5L//C2xP30nXWp6SpxXFkxtpR24kptIE
yRhm6/ADjB48dCdjX/PZiCh9pVdjzbQke/1p5e4jFoCepRu6i85TyvBkMILeXbVD
fOCwfO857L7gvINzWcxUY4S9y+WzoBwwQdlKazyjwUPWOP0SriO5VVjoGodqQDQJ
7UFgBYSidmyeBTnfMu78+P8CZX6NADRdwveOn3JIFzWx4cOdoWxy/AD3tRO6dT4R
ysMBtoqJomGzMVkecTYfMxqKwUFxfqY4benKD8ubsrOxy2bJ5XSzVm0uPShrtZH3
meDMBZGsFjDqJFK+Gd0YblfNBdAMsrXg8+5duWnBNJ8c2mEiauSSIbT9GRKldBt1
/payq3cKIvG6ChHPJ+6MPMtPdL7rnER+kql6pBPv3qGXXrpc/vNd3jiIDEUxmRj/
ZPx1tyD+VeXnIcCYhyBHnV9nE2GhpeP/9wpksp0XY4nu/10Bczcg+0dIm19jythv
hWggtJ75iscBGbVUCi/wPJblZxXs1lTASewmtjwBOEoVRhFR5VDRqSqyB0u4JoGV
puuGKmr7pW7siSaGTwOXZd9C5QhLhDsEK4Az7KzZSfV69MeQNw50P2wXxzia5tV7
keaOf9XrOcubA55vCrOtu/mx8wxXE94pSIyUn3XOk83xi/L8AHKZw5V2COfPBO70
/6gzDMJztfa6Diayt8HlFqrhdQXBiLTD3C6gFx2Xf1WF0b0OUBni38xNhmNVqycS
As0XM7Vmbx6XynugWnZjvTUcg/UcgEYb8VBC6igoiP39eEj3GSM6rEDJCFnpE+dT
2LftCV+q4e2DQw7vATGvslWvZChfoli89ciujC11dr0DVRm/+4KpGlTSY/e1tf1i
inlwBXJh0h9114AtOswTtDMyBRgUhAI4aIQW4P8fq9NkLRzQko8oaJWzILyTNOIj
1PrcAbfG8Z5sYIwY6lrT/JgOXyGwPyLnVPzizyfcnilMoIgT2mG/75J26tGqKDrz
s5f65dPX1xoeIUoCPXhv32RRX88ZTIeA3hS0e0EsiWeSufL1jrNu7tfCEnPdcWXm
dCtCfegVycjYZ5QeEmVxdDkhlYq4hCVMuwQwbuc2+rQ2n6i8MlCmMKw7IInsY9s9
wIbJY1KKBOmYo6zrfPKkt/lHeUXNpUiQqCxnB+dGZWYdXpuEVE5DyrlmW0m4mW4r
gTc1OsUajuaxCSsSqs6u6K1PPwLdbWByIF4ZglIKS3LBDPmwrpq35CF0HjU1zvHE
vFaLSODBgDgkfQ2QAz2QUGQh1hCTjYv1lID64vVUtpKRsFRL1AmOa6nwGPqznU4Z
EmVIp/upO1cnjlHzXNJEhjb9047GpkWG9l28yXxF1ZvzQ15Rvm8jZpM9NiiVgpUa
Pa5fTNbXSHnorRhCMfXFfUgzLcPjiXrG7VgLyBbkVcqTcsKT+JqqQJg7roiBwsT7
yjfoIAtZXCsQkCoPnvu7X5zFj8GIXcy2iE8mC+PW+5PefaOlSGviGSAR4Tg3EQtX
5ajy9tNFMXWYbNoNFEzW6jabP8oDv7hk/8q1NIbrCL3RfgEt+YOYNDRtPPvQqul+
DnC6iEifc/Qk1d2KXEj7SkjZlMq0MqLpOv7y47Xwwm9fYAA2BkZWuNKBDQVYJWR5
llOWdbwaLnyuNY6sOYpGmse34Dt0POYKUH7jsjcFjGJ/8IbA1QRhbuTSWGsJEN2I
NsKgBi2qq+WPBwJhm0MvfjwXYT1/ZrzccOvHiGtNxNltNC2WUbmVJgJe4AYKKhVF
1u9hUrc0p8C9wuxDI48WEmXcKvRr/F5Wf6DZhdE7oEPTZ0ivxQyEpk4TSnImYkuq
Zyurubb7xpLQjYGne2+k/DFyCFMxXUyRQ5I/agl8YCvgUU3nfE9iFQC/P8dmTze2
w5+Xns+RXNTiVBraqHyKrpVQsXh1yULRkkQS7c3dR6pIKqIGyW1l4pvIRzQds0kK
3+eB02e9b0OI/TZKVt+z/4EgDECMd4YEvgnOFSHuTs1DOSjOMs51YhSVbGCKGYbF
mZWrEHA3j9EiHxylIv3Z5aSGRdkbmZK4POa/M5vpYXWMXaGOThmO1urWv7Bsvxf/
K5g8Be0tbHEr24rRMeOEaKjideUF0H8DZmE3hyttW7VQQaklidGebPCpR5wEFRuH
S92irpX9jK8hDXiVrLZvNsnRatXuGX5L9g7Jp8YXs41N0YHernmYZUIvphPe0dEM
VVmrwX97TZbIdJCqrclxqbe1zGw6cVQt7L/lIzhFJZMxJfPku59gyuEla5NM3SrE
JHX5p9CO2qHF9griOuKCDuyS3Cqp7syIUJFRkHLBHcLbGRPP9vKoGMs6QA2TtFgK
Sf4Szri1dv2nGfxuYMla1gLop20OjcKMjovXG3FsQpLJP2eN67RjE7BJ11+yBbid
liZF0BPMw7zqD2HiSHBd6WKp9cw+S46Tijp/3ayujpGNjuP3giBFUMX1iTiXSu93
gcg0zUCqknzHPPxcSzcxLnPicxpxX8xbHe9+OIgxxMl4v3LL3TwbfFSDpc6VjL+F
oRZp3t/F4nNV3yCYym9WKBagYKQ4BoTtqo2TjsHV7ynoBiApLOGCjE5AQ5F1cAIp
OEQIFL/HAHrIdCIbeztkhA9VYJFedKNVSwnfNqsmUc4MUhNHm+Js9zGIjJJs51kR
V2CmWM5QSqmoRFuRp152IUa8x/M207Sh5xN8nrK1s0Qy7S+y207Qpv1PDTDaUIFY
sSVCBd5oVnW8WG/NFx2YLS6G8VW5YfaPMKOUBVnTrHd0E/QYMQZCtS7sAxV+AMn7
Ncq9g8pu7vPnnsKKR3Zt1iXpGIV/wipcKPKjjEmFFNkENTdBh5md+6bNqxzSzywO
fOPoDNd0FpiC8Wcs8wKLUqaXIBscoZhKC7juYQBPDYXZArh2vEBIphRaS1X0TCV2
iO59jI/4dbKUOEAjXU+bUtUcR5gNtpf8n2VfN+bAQDL9NxEK8Z/Rl1+GQcGVwLyV
XQH5VA6dSEicFgnE256+9z7mg3kd4HHB08iBbXXkHRDi/Nv7bOzmWKO7nP1H38By
ABZ/w3sfsHqpO+3/kbD83xv9IkQNHubcWve6xJ6HM6KgJkiDZFpTbSKBOtS4VjEx
fcwRx5PWLx8ejMiWYMc1VpWrgYWFyssJ+ZjrFqFwsXnnMzDNfTQ3RGLIsHoPLox/
9UHw6Qm4MONd9jPSzxiMbVi083zlj2oAy+1RPFES9EEQdOwEE+yuNzvEl/WbEOU1
vVdMosSOPfCfsoHKN3FTrEqGs7KFzytHRfKtUS0tiPJ+5woaonEkmjRTX3579vXd
+Kht2axqE6US4st4jrZhvCaeTk9x5KUmPJ9ELmqRKUCAtT/noTvZZAJ/6kAq0/vt
EuiG+StuCWZuVb160EIlCsqi01ln8cMVs99bPVXd8SnLgRAwDikyWspOe2TJE9Zi
j4GGaIJQpUxBpshI00Jk8Vq3NFG0zxWfdtRf2RmzvOhdvK+mdvo8z76yo6ELC0bB
91IC7lAS8Fv8e5Ss5hNeMFTaA5jTS4qtREI4ecnj0jO+YGWaQ2V95vc9u0gycYCk
nPeGAX1H+/YwLeqn6kS1VMatEJcvas2IBNLQFtgoADrE4ymMsvOYtGh67PSdAEOS
fjci89FslYZ+5/Ok2m2nWB2FSZvHrZC6hRfB3PLsl7qU4BZO5xL1eiAPb9GNwvAi
QnX3RoE6y5qLzzGPmAowSA4LMLECmh5jO6f2My3VfaeIg1XW8YFRzWTGGq5w5iV8
cnKKLk+NATUiCISNUcqolw==
`pragma protect end_protected
