`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PLZ7kpf7pBszuqdIr/OZJQQ+yfc16YAWTXAnFTVlMhzHv11rGEEmH2TdfvHiTrxy
grZ2ue03j+0FBI7ofESYLyxFvb1SnvZSH9Jlc9iq5QxE+506Ssv1KERp5+GSJ8rs
DAPbGQUfw+pFMgL5BYjjnKAOkRCfeV/ecdFv/C79YWHsTQsEoMslYvI6EqB4uJiC
wCmvKUGS840lopaYJEnxEdfwpRDcxdV0c3xjVntiaiHOg9YxHe8jwK3PM4yvvHrG
w1uEwh2BvI8OaMw8cij64qfEPm/mxpVd8tsqJQT0kz9Es97Gm9jXywZhy+ki3dnd
QJbpTzvcuS2aP175rDQqoA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
oOIb4eye4nFwQaAWp4IIpTeuc/gnPmkZLqZkIbEtUS6phvHVQt5DNnAsRUPNUsaH
T60eMVGJfCyZJb67V/zXSpK6OYHckIEB6w+UPo2LUDrv8mPLJ4S/PO4AMHXQLCN/
ADQcnOF3ioyZhumTlB1kPq3YgAGFtUDRtS1bHZReR4ETp5Iu7RVs1yWHq0Rl01v0
tDCf/CNYO70sNjsU7SRsy3JSBk4EVf9v4C58kxpjpvqGBRAlosRcPMgsg/hsn1nw
qgYqX5YczW2/CDEV5dJAiTtZiEFoI6+aYRpMPy7u8kLcrI6phkE3wuDtrFo1hRtB
2rNYCthuyZNaXRuiVdZ2tPc5hIJTHBSqiificEolTXCKbbsUfAaV9HRDpzcqUbYX
CtqWzMmgMCYH8g9okVg0WrZZvUivnDnvha9bBKtO40KOBkpPwJY1IkEqjAhtXd6l
gB99Cg0H/ZH+sMH1kUP9fwvjmsnmjbcrpw0PfiFT+nbFJwGNgLx1HhiQehxhS5CO
6k+g4M2+GlwkX5c/cACyElx20zoCKiUIOHq5lUlnPTuqFjigKVkajXP1EGWowHBc
8hKiNJ5sXGz1Pvbe48V4Ct1h20JNiGXfx5FGDPji7H7FrsTmNag7cc6RHamcdiMJ
ZucaQ6hAZu2i51qbNyDvXE0crLvsnlY5S8pvBVW2XjnOhemgT+LoH4DjQWTxXAsA
uxXOpRsOEzPNwYPYwG5F2mkMu5DDqG0gVDRFov894tUHyNF+KGLkR1Su2bs6rq+d
W38OwdEeoJbRHcEPaMKEoTpt+NP1Un4SeN4Vzee+1eBT3P1fBZBW/6weQnXO8g8o
/j5g7OjwEC4JBEUE2yrsjdCfvlezMmDBCWzhAPt7X5hihzzh9oH6kOzg0zW34Sl+
4Wy2NrPgasTI0oNsGBdxAAEVtyeTvLnAIewPXOXO2Zqrsk7pLeigWszHDhdFCCc1
rtyazEzV4FbXe4dBiLQd1xcL4koPkp8RvKTTxCqysltlWpU81OobRR1N2mFOmhtL
AoMKWmm+ZmBOYipfFIOl5SJuzB8B0zgOL9qM3mCcBaguuFUEdqTybYqEhK7dlfZ9
RjsoMc3YOQWjm2nyl8ThIzwhf9xMJ6rgrTy5+P/RTjNy4IduZCZNW+pWchjXHj95
ZKTZiV7uktHL+d6yYJRmgWlDcqz1P6Ky6GYouJfAaNFC+qhn0xq+0iZElwAYVMgF
6zQq1eL7mQxmKBVkS7rVSa/XB0rLFhuTSutYz8mPWX2+0dzZNpB8caUPsmjTDPTj
UivPPUbdLI+meUzxOhxajBunKMtvxT6ff3abk2CL9A155D7Xiu33Cgo4z//6SFlT
nm+/diP/DcWIuHgtSXYlbqVrOOeJ9PuAYW4YsvBOvQL5pxy6de/nLWcGfUB8bAZH
oZL2KZ6KA8RnnB9KJYV3tKUl1ami1tC3bVHOPbVeFKG6lkUj+0KLV+T54/SB4Cpv
7He95ybTjSqAK9Aq2Wlu/qwy++eVY8toajS+SWUzPEgEY5ziDIYQFqb8rOP+kL87
wvVZK7i9eFFoswlzhGD7U8nuAHUuxTukDn3QGj9Me4rWmOAathLTrkwa+lxL+B2n
MjBVGvmXPZH9ztD5qXlEJAda6sD9u9MlIQpPUv1m0JczLxitnz5BrOL+U13uP6Jx
cBpezOoeFk5pDWTKwtULHd+QBajvkZotk3+1wCFUFc0PTtTeO1qPUJBrysCPzX3I
wJ7OiV5lz7ROhV0JWJRG902F3ctJ1sVjhMDXAyY9A+1l+HxmC2Mfd6hkK2Zt427z
LlWUvl7EOVjRv9dQdnutbLDMQbStGG8fsnpBu87PB3iWQF34WPHnIyxZZSInrHvM
vmQyYbWzo2S5Nhgb1l36YOa2m5LcqUZB4Kh6fLGP3repgR8ugHJbqKMub5pqyQFV
HnT3Lp74KM6nR2licUieRQOOGB/tNf1h1cq02fa7Tl7p097F3nOxm5W3ai8BpJlO
7vvz6tYHm/yUFR4aqZxNa4Z79lzlDdLIad2m42l62cZkPpCNps6b6txInKQehhJd
NuIfqJTFm9rOdTUqoKxyUPa3C7UCkE8XxdY2V/RqNTfH4xESXbk/bm+kOq4kFvx0
FyLQqdWcXQMzRFEd4tvMLKiLj84ErlcP33/YiiQqTu5hxAAMmkTip3fpqmrPqcFg
Im9YIEg6oRaocWZlqKsjC8v0cqg6xS0nCNBxtU32MeYvzGFV04LEpV6nDa1jjQ9x
p/I9dDEHkPGbipKS6HB1y7Rl4TYeXQa8nF0/Cs23BXdVMsVija2Y8B6P2vGhcT/n
MEE7NcWJ9y1Q9n0OBiIWIDYSj2jsveC74BCx6BY59GzrR/mdJMnIHFGFvkbypmdr
hyKHMOE68Y2k3qBw9z0Q9MbdrWXSmDtYKj6/vo4ZTldjik+HyWckQCPbyqkoP4ah
U6g3WQBsu+K6OpIWMVOdjDzE76r9MPbRhtaCQ2i3BZ4C1KEq6qtThOB+ejgGEex2
zCvX+irRxa46NsgkjmjSCgUYTSDrFs/PYnKhFgIxlhRbTncShhbNiNspX6n6RWnb
0DtPVUzkK9V5q0x7TGmNlpxAFcRBexkaZER9AfU15B+2VolYCrUqo++ItM+1HLKu
lXJaAIDr58gX0phPKHG+VDTr6Gp0QZnwQZSK5kpb6WyEG5HSq57vRb41+wIcdynU
mzOg5Nop3IXE1vqiQeVPl3q7prDfajshPeosfv0KWZgyGxRAQSmppQsCHbJZjf8A
fJGbtZp0AkeD61O03DMpRMI+E8SrZtS5GyXqhmSGUIsI9B7NRr2TXqyu7Nt9jEMr
AoY1zicVRjYyeaGrOYJhcj9fjCntIBqXf6KP+gIlSNsSdMjKIHlFNfvKP+jabLmk
+EcbHK/AA0VyMnq/raIHLy9maiPCWH3VDiumUH6pAD1RFiSCyAqaDAbIKf+KTWDo
BItVuMwwG65QYwhd5RUoWVfmSMUmaohz6pk6mcqlc8gDfea138SZKx5kD4pGlzr/
uTB3CE/H2JoAuxGiU/8kFx8veJUf1yjAckGiYkdLP6B4h6lA+tCpcFNsQUzgCU5e
0TxoU1vSR2p3T2vl6tNahT8Y8NtQmxUA1DbgsxwCG0rjXSUQ7rTzdfS0h+jHX9zK
d9GL1rygz36eoqfksor3BQzn1JE7d16s6tmJLgG+EYmFqmQB71eHRpsBcqVyO1sC
MqKdlgEnAzjcmwjPhZ6Sx9LnZa6VdVjWpyPQ9ys9EkUI/Ekb4atXG+8siSv9VdFZ
L9glmINNW17z17bm9ynRsBk+agLFvkPy1AmqS1TUw914J+sMiMs2vKp2NYMrdEfQ
zBjbkxM6HLHIR6jM3u7JnyZsM5IgJzSTh272L1V7lw6T2guF1+sOkRe51qI8bHu4
6nrrMlOY9V3UVHUvAwLig1SBPX7qJhQfy59F02N0WWnh8wSAXklnEg2kB06cmwid
N+TIB3rG51XqY0YbjwxByH67hUxHTNi1jNW0rVwIA1vl13x+op9o7w8jVA+aghHS
RKCVZA2DgDNDpcejD5pCyWV/g1hVxtneGXPFd535j24qwD7/30o68ahup2mbILqd
OFVz3Yk8a90iEKIV2fto+Js+7Sf7AkMDtlI6898owJThB3a34v+lsGFq4EXkfNZs
rBAPwPx8O3SU7wwtRYtPdNHJAtXqFp59g9xwwZE0Deh/KIjB0sAE1TzkHEd9NsOQ
uFJAmQ3PYh3W6WQSQv2/acwSShVxCAWsd0xnFiYm0sALS2OaWz0ZiAhbq2tQ/6lp
GBID1D5gCqZbFJ7x8KzqlcDWtCFVd5ATZM9JkNvkCg3JzMQ0PWjN8Zn/x2bAdw+M
QN1MvlWocJHSUFpCfbUck1oFyI84/nISPhKkRp3V4uo=
`pragma protect end_protected
