`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KRZTx3/CrfqGz61Pl6xY6HT7Yu/07DFbNjN+VuCmFWhlRfT2OdcihVJvu7eGKQEI
nMfBAf8OMCm9fmvkpucq1cjTzgKvAKSHzdgMJq6X5RFMY1KZ/JpQG60Pbtv/x+aZ
n2kY/xX6Sy7VsshQmT3TNttBM2XTQsPJqnXAEb93HEHLGux53pzBSuQMgL9fbpdR
qMzCWOXmUjo1ZHS0w+9AXUwEISLnUUQueZTt0z5t6KjPIY3P6BwR/gZfv2H1jTnR
/vDCrk06GZhT1RWIGhF6lFVJaR0UYzByLMZpFlYa/P3VXgCihfSqNNPLT2ZL4LUH
WXwHH/6P/n8CFuA9bVz2lA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2496 )
`pragma protect data_block
q6KS21uncn2x0gySKXM/b45c2HQ8P1vyuz1FXdQezwJ31AnCz3LFOamdL8rcLhbh
t/zM6OCjuOD7Ve8+X+As2Vv+ysr1QptkOAcfX3zEMOpCyRBE5EsDkUQpYw77ZF9a
yeWBCLT8tCaTBLE3MkLGu1XBCq+y+xESMT9vATQZa565dbb7R75Vib9OnP627pkW
7nzaZxNG5fhi09hFQEDySsTK4rr6iYxYstBfdZkrJSFfSiXI0jC59lPM60db66Gk
SncMsuKDsjmGA6DmjD0v2Ti0/enzPmc781dm+ePPpQgqDkdJExn5tq03985Tb5Rr
JiVnIvT3nJdSe752SCv4MFgrxDFt6+IfGsvziIJyB7F2QkFG7wymVbC4QaY4BqVR
opTRE+rwqqTU8cSbO4n58YSTk1tdG8YfRSNXQgPzdojAIinBgOs9xEUhqN6EqmFV
NHd/gMtGLLC9EYGSkqpv0EiGljO0RPquhymKfkgl3k0T+bpgQuhnouSZN7LNhhHR
x+S1qW7EpuvE0cuIFCCZ6IRqZoYWe8HhS0K3M/YU6rqnjpdIgquaB778TLqbPWBj
3S7KpodBDe718lyVwMzMVj7u4ItoRKJ//zJIoYsJhosJdbaYo6pVXUq2bFy4pgZp
vFxcw4ZzPloI6yc1lHL6mtSBSfUV07EQ/WSgy5XFSEf+YaCtgQA/60ofGeNXCDdE
npvg7xaBJcqimaskbi+k0XJT+VBTaHDL3uQvmeX2KKIeZJ+LilzrpcZCC1N0Ni3e
AFAeeNI4KjauhE8i7JIFDSONcYxf0V6fZpYmOJg+NAJPlnjO+SHZ/LcKvt0cIvPJ
Ye7uan2vkPW8fHBT5vkQWjp2eW3ki6AOO45qD94yVQ+cgvWHrV6Mx5p/W8dbaU0c
y9+PbTXAE/NrL4i3fgLXVecikYpf9dp7dz+yT9A0anO155PwisdDXQfo46ZyLHjF
YXewgduYWsq8HH5QfZEEXTv7bp2+pjxtWxyWjjWzTckrzcZSCPE8K5Jx4EjeTi/w
CgfgQ1Xx+8wo35q+tzjcp9ktneJ+QHy4OZ7P5x85zfwKujx8hRdRU9ISKulqqL7s
cTAOsAUnZNeKQtZIWwsSHFfM0DsLicju2BW5nPIR1ZnPeRWYmsTTobfk/TgPMgWf
reOnRtSsK5cXZBlHvVjiOWqs8tVOWIWjyu/fTTmzq5fHdK+9P1BPnVTEVVid8LEO
8TZjNsJb2NsVwc9MrkscO48ivinwdTilh/uI0zSDTLN/kjXU2N7/HUyAiscEODVT
JUwM2C7sIyCI40zJavZLclktZ8vbz1D9/EWShSuZjn6pLal5DspQj+T7II1dC3hr
0s1Moebb4S2b44WymLbCPbbzQSo5en4llvPGGPRgWXoC/AU4MDMFxx63G5iPBbB7
L7knNPo1690uyGJ2vMp1GoMPSqVPyivHKVq0aUjUwxjd3gevpqoutsb9qLwbMu25
qIbJjoSY998apMSpkyNrYooAWedctqDR5RuyyiEEzl7AaIoIqzRE8jznmRK1FZ87
wqYqwDSrolHX+S/6vlYK71aT19wswbSO/4XPibI+WejWGoWNesk4eQX2lCBBzz4k
gWgy4NoUsjPVannR2QkNCkLSumtbQxYk97R9brkyWnWeAGibqWvqRlS7YfarBRyt
JD8jfMbuY1aMJl/pfJaNwyftDGMhy3CVIGrZeog3ma2JG64m4dZtyH/nMTyyNuKR
FFSDcHDsR0byT5f/8fuDyghRr4rSCOhDwml5Q3oROGoSrXqog5fu5nF54ABfw9Ft
CdaaEKjRNwnKxBFKu2HcWT2o5lmZyZHdMoyodSjyoOYjnmr0Pd0xDzFVAi9B1toV
/8T2HU5IS4+NRBDZgSFeAnEr6ZCnD/PTLIz9piPfK36vCUD773zZ3BpsbuKFDyw7
hdsaYsT7aArXOdHIRhboAKm8IgFhI4K3j4Ix9rl4lkFGsaG9Dg4DNzbWRjMg1Jah
L46tW0WPW43ASzkpARlzSPwDp8G3ve+v+s3huRxxr21wJqXyoaorqb3XDoC1BozR
6NOm1xg6ULRhz2wPldN4ASvufzIqc2excRR2qTw3Hy+jZe4P/8Oc8UaaRl/4vyfP
XZ3KcCPqxXOPFb2RXSIn6jAP0/BU/XGbl4EUB4ACm2uDHYdeK6w9Qa2Bp927kaSf
XOaHtPpCJmj5+3uIdvKc4JqaNxzV4w2hUb57WXKz3bCOkqJFtpWKVLTcvS/4ypTt
5KHTUUKWNsOF52nWa8koXqjGQutxkkgVCXW58Emc+q1AqqIUGBA1UOTisBViltbk
BymS3EfSeFDWDlK+8TLXtdYmThNnit/tts+7Mpw55fZwy7I4L2zzA0QBkfEXPpY5
apGYojqGi+uHIza0f6n2fAU+dIgtE3kODAivmXxmNUBUr/5GS6ohpQy+Hq+0e+Gd
NlpDXTQJKwKb9Lg1YPK2Hed5b5KqzAVz2GB2BO++A4pKhR2H+rbv895/WeGgLxgn
bZ4YIjRnrQz/b3mQOn5GN94vghYHkVO7kivJawcMzyrqAQXYbuDYdoHY7j9ViAJ2
dE9OUyuCZ7L4d/dU/tHdR7ep7vpZMxjZtQVLwhss4KOEVF+ff/F6DhJ0QhJ3jR4h
aICGm3LhOhZqqrJSPlfy4mJagK/5MtcPdz+S320pnfx4BIhWQRLArHn88sqOFqD+
KeQiBKy7HBPKBSUBlFn7iqX/17GLfBFnCbYwTGD/ZwYO8+NSOO6ye4vrEuDc3mv3
NJY/BaVOe/gh/g9+AfXy/dW9IwAMaIvnis+9Oj/h79MIFajxiYrYnydtYqEeJaQx
gXqcSLF7zQYtQtAjKM98+8p1VaQg8BqSESYCbSUoGNQma4Ton91nWwBXuvej2peR
RnwSoZKpEDUpkGg0UR1gz11PKJcrSCNNAW34cxqfaW7MxBvUZY8b9g+isNJnNDW3
jcCxFYUYktqVLKkSH7oW46tTi3R/PHb9hhXj1pKqItTLWIYQ4ZXDpUieK0DT1ZW9
2kdlKAKTBvUSsk8baPNyHhbU8NfB7eofIeXlAXPYjtGjiY66WrqVGYLgv8eqUQIm
NIdhnAB1cF31AqWCHHxyQbb5SDwT0/Id89oL+82Ws2ymeihzBE7HqF3HiFxc0jq5
GaGK1xJ2UjTvVxXlwVsR0nANIMykNxnDQbHyh8caIhCUQ3R+k3EghWUWGJTZqNIa
TcrxQRKKxlYskJRpZaR8EnS8sK/pPOQTNZNyzvY7KVbO/VteVhkYUZbQIbhcWp2f
makl8kFCW8PCxS/8pzOPd6X+LVgw1UCSlhLVI7kaXZGwroDFpBHnT6IL1Z84Hqpk
`pragma protect end_protected
