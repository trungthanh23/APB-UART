`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
s2sas9riRcLHdpPQl/rmfnGL5EzxS/i1GDVg/INfNJzc4Jvf+qgr7AcxkWoF61Uh
iEqd609lLH5ErAAaLE2myajfuP8DMGaqoduK9sjCy4ZIKtxTvm01ZZS2GJ+bMnu4
cuH5EOHuu0wnh6I/Hx7hhrweDhkvCzxV3wZYxv8I3Sudu5ZwwGTivwSgmS37i2ND
ngMbDNkIqJdB+hXcPNYShOw8rgCwOkYvWfs/7SnfuZbv3YK0gJaWadm18CNMvmVP
Ll4TzcucmvLTM1PnV3z4WPrMWQm99tKsLNplORAy2aAZudBSr9otyn3tQmbiDo6t
swek2uTrhTvkxlT4/MuoXA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3360 )
`pragma protect data_block
o7T+fBzQhH5pnIny8jRTjw9NO1RFj1jDGYPluIPnAuiHsA+hcRzVZVvviZQSdnI6
meIiZXmPk5BCLd4ELBX22fqGG7X4QG7kLwUPgFZBuhI/LI/ZO3zyzLv08Ow6K2to
S7eq4d+UXgFUuvYLfrbq0x0fzG7+gwhrWgTF+/5fYy+hMKC85qrx8h15BhMamwGz
9zfLPen9PcVLi8o5G32fTUc3OQhhJ21VltAhMx/5GCupbH6J/1xezvZI2e2WulFa
4UWaS1C8fhCbu4Wsdads1mE4OqnwdQ+/SZFxF3HqKiTWiK05qXdN2YnpdZjZrVZm
saq4RI04XI8rapNNkcMytBkFYJouT+vJyy+Hpnv7lhrUc5GagEP8nnEoXNepZ309
ttGH/nXQUJKrN1D1E+4+PnGxk3RkaT0XNIEahYosxuS/KcIkcTjVIbZiJi3iuwlS
XK+NBKNz5lpZzK0lAxfOgtUnZlEfmgAwEQGWFgiE3pNisMiRLktgsc4ygA8O/M0q
YC9RuxIrsFgJyIvbJpt5iuzKltklPByMc7D474WCf78zteqKtHfFSUZOqnOLGpST
LV2raFbhiiOPCAZw6tONrja+OikN8yfiN/d4PkF87oq6NsUP+0VINotzMnzNu7Jw
2VzES5ZNbyLrTrmNB61vG8BOtgv8TeR9YJQbf3576Ug+poZuCaIZ1bcJM0FEhZRA
lfmn57C72Sa1qyQobsD2psO3MvIQPnSP7mabLWwUJSRMJWRokzh5aeKQQs8Vytw6
3K4PJlQKWGGMUJLaHamJaci8JuXscxC4B5fx45oDnodOHtgrfuFXZ0q7bQsaXq4b
TLG4wFy+V4PpabqNjUl0mQfy253xIHl5MUDxxhBiUgtuYJILUCItK/0u+ql4+RWL
Xy31x4w6IujkzbMHNYT6wKAESmVQ/0vByMePPT7yUQe+4E5kPugvC9EkJCswQXdf
/mLnWEid6gBuT6aZVbeJ4yBEf7oP9Xqp4ZPG7AHkyW3hT00PsYP7pkRVTcS9YDxW
ZdCokV0ep/CYuL6i/wn9yRe5XrUVVeKe6Gj6OeU0pdbWFQ4Yzy75N3ccDz+NMqvo
3LthvxT27TuQmKO4HFiTat9Y8Gw09YILd9mGd4L3YSZDZ9qj8ghSGFlIWphFhz/7
591211deap3TeTfzvDcWAHsVuebzOU+ZNPdvL6t3nCEsTEYgclEXN+kH9caItOd8
QktQ7fgJfogp+rW9G6FxTjudlwsugWLL56KikUVQ/Mqqc90lGpKBgJv3DMEK5IXH
LpfqfPYCnHBPBW3q8UfuAj3YHxBHpPdi+z0AdVWNtjBLryEROvG9zhDd3rfwiiZK
vASaswubEg7in44I84VYQ6LOYwXVKHtIzljYdeSQ9NoVrm6J6knAMfD0QEOXTGg6
WobXJmef5FQ06pOos2KFu8lx0a3hL7yAzjTDZGgSly8zZOYQhGbaojU7txOPSYdN
+T7vT0n0j4umI1l0j3xnKuywUuSZql+LxQTmmcK9RxcpLx36424ggACbvplzcjuZ
zTLMJw8yFYjNFbf9tfXucf3UX0uVkhYcoJJ8YkjEdKdud8AYiqvysCqEcMCjUFsm
+6fFW+FLqyKDc8kD3tk8bhEtGy4ljT5ZBfnHD9BCKA1D2VCdP1Hekx2D6ear5RA/
QdXXa+Kj2nV+nRVA3x4ezHKebErBf05g32bRrvnHZ23bUBfiLOWBTLTvhqORDcrq
bfsaeEIKrpi6Z/liSiDS1G7fHHqrUmU+7uxCiAu65XopvKpd1im300so8dFEn34o
CAjSD3PZOmsGv9EL4RUx/2Lmfuu97YycAO5ybqbrJT72rzjb9ISZSsSnmrPsZd5J
W4kNW7LhhG8D9K5IzuSB7za6PCn1YzSJdDdPlqo8IC3qNoRvcppV1ynVD7AYw2NX
3NUAOAK2ecQPwesUZcw2GrDOMjcQHRNdWco4FeeYm9e3nq6TTNCygyUx2o/92s6U
fF6fmdbH66IABJCAQUYk3W6GtCL1Ebh8tNiO8/dNiMVrY+MpYS1Rr5uORpHLxDPB
UVn/5lQw1CdkRBQwfb1pE0nVOPLNgcs+IJJPexOjRg5CCc8hBDzNvgN5aj/sA2iG
6Jd6fTtomVtdayUN6IKec4mqzECahWwcSlWT6i3FfxP7LZmD/gok7hbDISLGTIoN
IUD6vK9L2r5xNwAy93GdzbxyrlQ8SzdrYgARtQDYRGvb42P2lkqcOliWYW6Z7EXh
HBRmOEPdF+tHAQxL9iHzwLUs3+gZ5RLCtiPjh0CXWszD7Xim2OHV6SViD0yOPqW8
lbh+7FzZCzLT6fWBX2+rc1br9IbCLEcPcGrLIFTfqC43keAGn7ndfaC30D5lqAyS
teZric0XvKLBeipt4gbnRd5UK0n3aaj0cAiollXUjHdg0krn8Fh8E5o5as5WB6H4
SZ8CayyhWZqBrM3ZG133dGWN2VESLnyg+z4l4A+AMgB8ockoeLDc3iSE/uyHnhMk
znuYOhwAmiuUggkBZo+sagq1AU3ifqMpTOZuhvtb2VItmSp6gVYZepi24jrhcMo9
/HbyeF9d+Xxhao0c/BQ+ldwHkeAwSkp23EPEVHUIn2PlDWI3HA3EawFQ80X4+nRS
hn67vZiD7WLfAJwjVtX2ExJlFxHrNt6jPs6ZOK42lhPpqtO7iTTobO+V6ODWuy8p
P7v1eowzHHBSHFv3Yo1UdZjd//gGEkOMNrhTS/1gYzmVATTEa0daAGLSpQIlTiWp
jKmdr71OoJZEG63Ft4fNxUSdjJZUYqzQI3fhmPvJTqbfWCsgJ+234yxXZ8XT+c1u
LEoTPKG9NTwwm4UjGIssmgmgSU2kS4Zql18KLJfuF0GHHZS1JkQlo/nUHymbTVBa
G/SAMdqKkrs28KLEiKPnDJvWWMKnke5bweVcHNA9o1lmSLf2XxLO7XHC5WBGS8iL
n3OlbTQ99JevP3O+BF25dZGNMT92PvjR/QctuzzD7VSMhdhV9RgdJDSxZmZJM9tI
BwZfzEd0OkeBMv4iPQJXDxKUIO5fNfCxv6M+qtpAE2YTZqnAvEMO6yZoBWDLcMr4
QgHw0j/Gf1gSrU9PZdHml5hph7NUP8xlpZkSI7eBWLDdAAIrf2G+hbges9M+bFif
8R9BPMznbYerxx2wZsFgGPToNn5N1a87K5TVgMpuxDdenY+8oemm0o9BWfBIZZXb
WZv1v6MiGKbfeZiK+anrpoYygD0dhn+ZnCdcChq5bBOypnolWMEQQwJryjHW3viQ
UrhlPuaZ62Csou5ZifEm4byV7RtnuSZP7a5CkGjlu0SBBoIXLxvEzx7CPDcMo7NX
e9460rP6LbuHW1KhoJx9x0EEAXRDW9s2W/WUzPnsygzlKL0C+UhTzCTad/XEA2ss
7CTBkpP2QZySLaIEW6S5spLmCWciuY95hTmoTzKQNxwLZaRdxO1vtOipSizppoeO
96dPnwS/1MTvCj0DJhNWtDIIZxY7wqAfijJOiqngapWeEJ/dwj4Pm/FsmvXlXvNS
6PLVzKur+SqHPqvJXN9oDH/sLnZNvlZhlvoJ5Z/gp8823gs9uDHycKop2kEHckCU
ai2v6zCQNoB+b9ZeP59xHYt1pgyQfOTqguvfCeiws1AUEzPnq/lRQrTQhmOVmYED
pQb2pn17t+YLJJzPn4KOJKQu4EA+ww1OXS0GYv1bBz5S+4q65Z4gLNrW77ahe/8G
824P/hEg46FnfyU24Tyjeoks9DOO5S+twWzg9pASuidrMlZjkn+fs2RCIXpI/ppc
x5ubdMJk0Qa7Wj0YvNC7fxLCCcGJPvkHNXUWRmK2Ql/Xpc3pTroKI8BCJu/Mlk2o
wKy8FNt45CtTkqSq8d6kxOueH3woIeGq2C3Dp1lWQQBpSMnvZxpuPbqMsQK5eRLq
IjCd67zLZBvwE+jv4n/UOqDKO+RlYW30tHUQP8Uw9aYlmzQkxe1DuHKucnvZZEVJ
Z6Jah56wtpO3n8dz5wt+Ylf79zZmQHk16pIzBtpVbZ6A7p1l91Uk0mxprMZVkZxF
5nAI83vXRrHs4vplq0n3KS/ueLkMvmGQfOVhIuqYqsk9BbIUe3gsBPu3SNDxNNVN
IWv84N5fT/D3u1S4mBzQCQBGiYURyYXElZjttjeUdHozKbUMGa8YDit4EOGvngZA
WN3wyAj8gKIU/v+R2W0YVc1uSqnc26SJsv+F6yf7L1uHhdp54vNzVajI9H/oPDS0
4hAPMpJOnslEM3BTB2im4kvOPH16EmyHB3FEkrhtQOTXtraFUzd6d4KofSgAlil4
BItQOL6C32y1rFNbtqFmkPsSBogp9xravk0Gble1dvAdrf8VO2H9v5HT0kHm7XQh
xU9XHy/6LtJfsgmJzKTXmOSoK5ZAVICzuqVhlcISW4/C6WFQqfHsuDW7NXDPTMNv
iHhqzweKUsGgY4n6bd0qmiIrdjiICCwXtaXnOkKrhHbCKuflzhYel3Fk2LaZf+Tb
`pragma protect end_protected
