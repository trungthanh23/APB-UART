`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VwMYCtWX/IZYWchaK6jdiU678OdfwDrjIZGiCFLCpmnmvICf68YhknXyEdBm2ISt
FRcKeb5XkH2B4GkMyXgvHvj/TNap+NdCfEPnwZCrcnIeTSHq5gZkOeEZ0/2t3xBR
l3jhigx+rn4SiDUgK4ObpQeRqYU+vIWumAQQf7Pd6ZYLSzWS7XUsP9yKaYO4JHsc
otoXwmzSu/68a2obsUA3FXfY2EqHb6Mrjp7VuvzR3YwB0hYynOFUwK8IOS5DiRNC
ATR9F0m/TThrG2h/qe2kXvCUNNuV8VrmjgYyUcP9tRufeMHs/BHuu2K8D/dVYfuP
byEVENO5Hu2LzAY5Ugougw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6448 )
`pragma protect data_block
vU8k6Ebck0AQhQbv2i3DSGDwLMBEgYLuNOcdNPXpa7FBdzs67MNUtdmmWrnD/E0S
NdgEPZ8iticAWWt1UI4ShN7ZbK+xpC9tTklrdEgXeg3uRjcOqzYKtiTVG9kh5gAM
kU4cBF8Hn5UemRQu2/pDniUt4O2FlZaQNmgFEpFtsmw+Sa/0VbNBQVKh0gggQ6Ef
9IX0XnyOln2TGA+HpHz/Jpz2uDYH91EY937O7TisH5IplLEfwZCozrTAgMVPuc7w
9O7hBTotxn0yaizxP+XHBXiE91CeGvbDX07BD0T0oXEahKKqWArlVXTLy7YZw5YZ
5ptpdY2Ffs5jPymEzs8nvM46ojxiuTqunEi4j78SyXmz+IkQxE8GWlu2q2oplq9w
bfpAV4MgSt7auWXZ/jk+6yi7Q94Zq38Um7422be6LFnGYEq+Aic4QEm7gIzS4Sem
+BWZyuP8FyLuyFHR3ZR+at0HMwddB/9E2xnZWtZEUduY/ndXAxj0L/q/7ljaCH52
/unV/UnJCgKGnyp39H0QnN+15VJJGuJEkBRHsSmHmR/pHqfVTHaD0RaaMCqSo+kk
2H0DxdQIKpL2Zg3QFZQocNldRwNQE/FBobi9GEKUf5EJFDUjmTMURnH+vN1ihFYd
RjsynWPXAzTcNQxA2GKwic+j4a3wTSxlKn+ZUh4mAq7YmYcdy84zjFjMDulgigiU
tAaSkb1h9raXNhdw7EqwHcj7XyU43Rpq+6RoS9vzJHedQ09L1SgfCqeZ1B4RVLbd
kI5+b3yrISxbOnR6d08aBbMrs/U7TNC9KLb+vnKuarWMxoDfQW6sjMfVVqZ7h9ci
iUteq+spJ6jSq7o2COcMhRAljIZbrkHcr50cKb8n5gM9sGPj9zFxr6FYXvU0UQNj
4OF4s/nvFsJvmQBINjpFPF8DimgzQMF4uyT335DI/5b9s2xz15BdloZhucsloI0l
6xzuM7XxCCT2pT8Ei4H/qeg8m6VzhcvxWNBimCVBcC3YkGG2uYj/mqYHdXauvOAT
yPRhXvXMvUlZEvT/LHEOUq7DMu7z17WK0MO8vm5nhNxHDDKdcc12ksnemKab/+Wm
0ntqvdR1u9yjrj5X/ENEnImUuqOpQVJZp/UsD2t13Ed2xe8X3r0o6jTtxgO9K4K4
etb5qtGyQfjbrE7EKIX7VDSJAHXxucKKqjGH+u0GOzps3yaT+I01wnta3w6VYKDF
ZBe1CnOf8Ann0K6HovRAF53C2OxnSHAaWrQ3PaHeIBkDIKaGN+7Rh02JU9E+orzd
ILsOXbK/Z2ed/1FEa+edL1Sp0sCh8CifuGNJsnSv/xguM+dKrRsDWnN/pVBzMbMK
mJxP0O73aW4TPMKnW5tJO9GRSRPFH1REJUnZJizI53jNs0eYd90iaKCWFI1uPFMw
R/IE/F6f+JMEt1m1e8tqFz9eIvUktcEsju3ObrLOceduZJHMdgcw+k+rvpwAr7Lb
nx7RMxoP5kr5eidZNk7nKTRqz3Dm/hWLxV0xUgjO7IN9V0QQcEpbgEnW8dy9JwZz
rJPa/fGChp/SIyGwEXpdo/pbSgAPAhXKgdHUS1xQQBN2W2UV45FoydYjgZAAvBG8
mg+4L+KAUE2QntWm0M4Zj/z0K/QHQIHrkZHnL+ivrMXoAWgaw6PwQolF8MlPUbND
YyUqMTLDbJAC1YYbHsQkO3wOgffJe0OiABephWcGRYV3RYwHJRZ8cAI0Xz2/LFdI
pgLSamX8RJnet9BgJ868It+aDaSzPb6stYEMTlQM2jBSIOepcPuXo8iVZ7q/4PDI
M3EF2JnjzYJMKM9+4FWXms0w3aNUYzSkZetkfKt2lwTYW9fogLUZl9dPh8p5gshC
TfN9r8mzM2HGRD5t1ITRchCCvsdPc4CzjTyAmIY0gbBVy7DVemZnnCy+9qoMPyo7
/5GpmpQFIZSOJ2q7c5pJH06LZ3kthOd7z3NlzFMGPQSn9ZzaFsZ2jgiE+ZWUviXM
OVvliJiyvJBhxip58JHk88p/xffNHnbuKzY5QUEUPmpyXU0I1fhTGbMyUo4LAO9n
ZEcfkKtnO757xhTv6ssGZTXd3HGgTXpwYLt2MHfmBKA40ux1wnlkj+UFqrvxmFlf
NUFP+MaiDJALpZnxJa6Z90H1bC0C418MSuezINvFSFEckHtlaiaTrYJubX5dIMtS
uIjI/3Cu6FIa2G1CHqmiQQdLgxIL8hXp6xc2xsQ4P/QlL87QdxtSntiisqFbx2KH
Ve9ZUkWvlPk/wjmdXNgyK20o4HnVhKftibPCNH6MP6Kn5G1/0Fs5B0TthvjrxInM
kgop2/sEFoBmKMbVRaIrZtKA/tFWckJCg+z1KXHCPaOf75k0g+PWUoeEQz4exavP
lSJqHf29J4ktDiPPejqPI117j7SDh6NINTgcXJn7aAyBw47A5lq510uc/3HTGHbB
/UgWehObPuap9/JeKzFzYI/mOYdGIbP4i3BrDoW+PiUrenG5UoIqdIUMuIP3urTi
/angGBGiWUN1hNWgRWCFPXZigq4SjRaTS5pcRurp/0BkSdsd1MQYFtu4U7v6xwvP
OhXk6Ykwstcfni3FvpgUOpL3ADAJvSm+0ns++jruwVZ4DMFx2R+MkHsgp4Q39JDL
6SymuEu2tKc8v28g9Y4vHbgEb1ioHeCLOVs7WQcYZL0fw48ChgoN1hqc4fUw7BWw
nTY/+6mfVBCZdFuCtKxh6T1Qm4sRrQ9ezLLn2YPGlbbSguthcgEqxFrSQJidWRZ9
26nv1bFb5a7Vs/M/xwYLbM/0WlBXlkp0JeEgK8GGhDOgys8bNgPLvho1BW05lX/B
KW73v0ymtlumN6BumY1PyNpq5ADXirj4vMNCHeaVJ+KbxwBa6H1WPqNpUjesH+Zq
VOvqZY9ITQcio5X6nWozD5ivhBcoFBDZIyEe6hXq39+WZ991S4d3T6SW7aIE8q2e
5dE4/L7qVDChs8Haz3nJxWiPWDr8pBXOhv2JeDQnfm63guh4FQ8r7+zcw5cdnNv5
Hj+3AOAXyl0HVfQ+YQYn3aQQ9Cfu9h9d7C9k3+5Y95W6WEouUFjd9nn1zcnPt5Zz
uKxRi8vh0BBbGrzOknBbTah2ZFY3RNFQWXI6ihQx6BtnXfQu/BtUKPyH73QZg/Rc
BpYSNwTOqBUqjVbWOza1HWKej+TCRDBGdwn5Pg0PBjqo6b3zqR6M7Em2YShija+M
TFEGdfA88PqW/SlMEwCYr5CO9C+2g0lQhe1Wtkm9rHYnN4ei6+mOF8L8cJiUlazd
s//JlTV4YS/E7SQw9UvOGDw0f+E10l49LjrZWluhjjipGLk7h73KkrkIKYSNj24d
1GR17aj/g/6ZQIon5FReNztmxpT33JOpDOliMvW1a6Ebk39I3iVbDfTkMjP1TBc/
lNjWz55Ip3iN1SxVHl1nIUeLvJFQNzU2hz534/YMIoTPlCWjhyRUtS3nWiVRRDTh
X0gNmhwqq80Zkce0+dH90omovRml+JzrVicW7fA+9vnKRMtPDGtD/nZQKJoai1xd
SDIkeaYULr1EKVzoaYyMzgMBxp3kcHkGic8ny0j6ja0qdrlByQIYvrc/+iD6R5A2
2rz1/9dK8VhsYMerzb5O9VFX6W6oaAl0Fb6RXdM0ZpjnDOCkQnjywijbPGbvXvos
d0FQNVr7WvyWyAnLCzmJ+G8I+UjIpyr9nT8p5riVgYSB8so51Z2QUQLHHGHveSGK
q0mJsRmd4OpH7DeS9AkF4jrIp9OO/AIThlnikIY68SbyeB4Q7XnGAvo6079vg15m
Hf2/ii7gLySe3L6hLqjp/YtPM3+/S8aotu9PnyZY9P/nnOhjoAbHbp1BLyiU7uRs
ztgNblnTrcy6NN2ptgQK4JbJQLZHIyXpWm0bFnbfsW088W2unrlXcJkwXPbAFPKr
917V525Vzyp4oaHsOtyxNnQlVCx5m+clzbXm9noCbvCe1AaCu+P1C5Ds1qhD8EPU
0Dx16P6hLLu2IaG+Uz1eJ21hWA74ilr5BQRS2ujdxD/ADEfE9fXLWFuQoyuyJPt/
gdFPod4qBRhvjzF9nt68p3v+hfE1EUIiDg0pWHvLkW1pVYroAGV5KoYSZYhwd7oY
4Corn+TioIX/mSqX5XQJ7q53rXFRPRVnV60/95v4563pTMpr/0R7YhXWT2CDJBWM
Ac4lMkdXroiMPUonITAqWREoWghpXP+2sHznBBuCrA9pEbDhgE89oV9vuz0YPfnj
2d0yithUEEAtCEuymfX0QaG2cAOS40Izy3Q1HHegVTMv2Zux8wtExL9VmrorGGdw
lCH5ZlfAsNryHMzrSMg8/D0F98WfFMPP/aG5HVgWGcwNHyFhoPkTTvRMwQx+ljlz
cGSBTU/BQtMTrqvqQnamyAj31IoXbdofmfpKMpy49S1iQUgKy+LexXo7ZjoM4xvO
/YAqj1ucqvyB8BOrt4CShl6gu9c9NTUloaDskvYQu0etjVQmxkiSWYpqcHbQ/Q8r
70S5Z59/3yns3Xo20CqOIaenITVibfk/L3cMnW80Y36/4DdGQQoGkjKv5JC6RO9q
laM8myVSHOxYzEuxgeUvb543Blod3EMHi/nx5ujRxAabDDz5wse6f4ikA2qt6Lbq
8dXER2pfJvemKOckAwZ7SF9luMsWPTWIEGDHxwIl6pXJdEgR3WJ+9/SXzfIv5Yim
wv/hyPL056mMjJ08BbsdA4zRo0+3Q4I9c3qBAzAuBylf0lzHrCl0B5SlD3jmuHTV
Iuuq517Viu3bizEJ1okcGaK9CCbu73iyA/X6upOZlMUV59dk1na3kbg9Lu1YGWMb
/+RdJyLdl+qM2zrIw1Mf5nvyj4TAfJdlJ1xB7u39gwTQK6vGyHPMZxfP04tiry4R
lW4hvE9v+HCfzNq3hTrF+5L5EzKJgDfIguWh/6IBqgabdfHK13YGtvSCgW8YnzlR
IXXdKNWkqI7Iowm1iGn4iRC0KDhV/vW3ddu+IeXGwGFTV+4QMgpgMNkISFICHsaY
99fD2Jhq7gbOWRra7HtN6mN1vfU1pNj9CGeaA0teRimpcNpJKspyOUKGp1VI5JRu
8Yacpq9buLSaxAhCMYto08wSlMPBJ6NnMwpuRIDMdM/Fvne4YYWa3FMCWT7G/qRx
FNyo0a78XTN9txz4JGUcJozCSG5GCVhV1ZFQvt5eqX/1Y/Z6Ys7AHyA0ZTgDSBNX
4jguHuO0B6Eq4uGXewj7imSFXd2T/XZ0M/qmhU4pK1+nabL2a7x/jet72kKOPS92
w6mMubNpSO6lViiKWSlxUWawaZuXJACsiuDn3AIZ24mEzTXbNk96GnLA5XRuindN
5HAjxwhoAjxs6Jo53gjXO4vDPBXhP5Hh6rxEkJYznt/G8ASoI4EuT61lTGqQPagC
gbc3ZhXxpJ+1yDxVmc38Zqf064Ewy4o1DvGwl4PeI5b1GYp7h+GeXJtDAGIxUBEE
9YGWhwK5Wl/ylGypw7tpmPZkvkYopqYqIwWCX4mjG5c+bAmuoBkqt8SMOmBd98/g
QGSWs8g950nVFYaMfj5w/4aoeG8hnCln3oXb8jjWnUz5XQ8Huf1bLZK0fObzc919
YyzojEvfSItNbLgu9gRSKHSKjXGnNyKBKSTDkAveGNMTm/deMAVRIt4CNkBzcizW
11mXOiVpsanwpSJHVXXi79VC4P1smHe6lwP/yr4dUl1WVNlHfzWF2KGkjaL+lb2P
sofPLkQGn2+wbEWBuWm7FAMOTnBhzDqd/t3JaOCUQHg22qMVAAjI6yHFn2hWC9DE
yWnLZPoqRhKFA22wPhQSNdIaLKgvchxDbeQCa+v3ueNNZ2ikXgTlmeLHgiBYvTMl
tiDSc4F810Tj7dSeROcj4qkYFhm4t2MrS6l9cajOhp1zHmsp80gEColOjtrKJCrh
36bGPE5Qilu0yyzmdBTFLp8G3s/Q3dewD312m1gYEvniKxdhvQt4OXLiyESrpFej
aAzorG1uzBhKZQI2+bv9R/Tmk5qOZ+K1k8clxLep/+/hgee5pOYqpk0ILBI1OyVt
XpFEluBRk3wCrY9bZLNNXgJFhgUE2djIF1pSc555FI9/kc2VbjYc7NogLyg5N0HG
zktP+Rnx5z/q0DYsiBufs6QcRObSTRdKLDnxAWuqI5rsHzydC0GYtFyyt+FIkIDM
Cn+3+hz3bNRAMHzk/9/ZnXYhVBjjdivOJ3Q8a17TiSQmiKfBeS0/YAMk8ebKDubL
UfFbbAW55zB2cjAfazawppMcT4UD0nas3z+7trZuLi7za3auzTiC4Z2fvxEjORlb
hRFfI4731+4hgm0cLvuV3w8AUlASq8EagxUUnymGYoLhSoTXMztBOjL+nXssUs+M
KlXf38j7bqIpMR1ct4ssdBaLnAhDpVFkkVm56l6gIpe3Qd/zgjHhno7lW3F9vyyL
EayPtl+lOGju/aQShXghubLQXhTkrT2E1YWLJj8Uj8V85POhg9CcABBMlRM3Bjwm
pNC4kA01p5/gGpe5xKg5mmga1/Bjm8tZcexFjxNct4EEt5xIZzihNLMQ3k4r44Pl
dYlJ/lkAcZGLv1kyy/xIWGF33xheD+q0ZJwZYwj9uYhSxq0imisRtmpM02i/bgWR
b7mLhdhQ0cN9QcInwXISJpiGuL+j2EMV/7MblbT2iBObxfEUMHrkk0IRwnsN5A44
lf6MlLfzXUwB+WaHFP0PA4wm5oiZ7d34VG1RkSv1dJ8AhY0mBt0nrSKfgreA0ZWK
xPegxOUkqPLZ81ped95Y5d682o6ek+p7zukZ6FyQSun6DS/10p35oAGWZGGkz/xp
yqk3q1QcRkTCoidVlt5UAtFY53F8IQEfK0rHzMQ8oS1J9lx7jo76zbmro9tE++AR
rTLyGrrgL5gDMmN+kSsjA43vgXclzHW9RkMuqYug5ougnlhudBPYwrwhxReAVjEL
tJvuYqX1bqB2MbBqe2t9qDGfTgll4MwCRHFwqjIhWHla+6q17RRV+NtVH6rXPH4D
NCueZQ6JN11jNQUynqjRTVSyJPgfmmYTn2dXyRl+lz1+fjmCbqY08pKVB/kI+ZXH
0Pw1oqdSQf7ME1eBErWLLqkhv0BgXyxoel+W7MNbK3xCF7JfyCosJYMl2eVietAc
rL8i7+uBrxCo50RWZBI/qi0inAdTir3KB8TDAdT5fB4A1TBZin11T30Cn5b/gtDA
7m9/vUKkv0G5xouAM7qTtvfdsVnZcV/THziX9zROdoaDcG4zFKDg5p75869cZzS6
yRxZ802tSGCz4xlKbdxmRjdKx8eytZODAE3B1DAWA6g4V7S4711t8EFrkS9nus4X
3pkctR0+ZW8keUXzt8Vm0rD71B/RVxqYkwBy8sR46VcFmJOU6kCQveT07i5NF1Bp
1xjUMnoGjwE+DfJ7h1DH5/7+uqTLWcyag0O0nxIKBau8Jgxur/Mc+rwMLex2K7/O
EqhCknCMhhxYNlXoIgJ+f/P7Zaq9p0ueFgUtnvMKLgYkewaY1fByfBlNira0Wb1U
ZWTnrZXdo4soSaBazqnCTubaz0dBDHwNIpX4AQHLjTDNTEndHK0uW2H8t6As0uth
AHI7F7q4+ptsnC8kkhJZRSUZcAx0xtl0dCtqM20aBNDpmrmYmt8dsB4O03fAAny0
XwZyX36v6/IOEGzkFW7bIDBuNInRu0oOEPuZDGaTugu1JwN9CTz0cXdTQNp8xrIm
6RvQi/lA9zGx+lYkG0MXEg0VszDSYPQFg71mYMgdcTdX2SeC21XhqpA2kYc5GjRu
gA7D6Z82owwAPI704q0dj/UBPiY9+VbLDsaS+0tCQC4WNjhTe5xNTNqNU48sKdWY
uOEl75Smcm9ex1owN864byq5YvIqGto3rxfBX7n5sY2WH4TPmCVtxR90Ko4LOJUG
nBkvcgijRbVUFZLBWQhpchLHPHBSASCO9SwRXJ/JKN2+JR52ZWqezljLQXvwt9cV
FzhTt6LEFotAsHhT5JZKNX0TmUy+mdPHruoS+gyTv0RiuE1TdTikNzo7O3SyaShN
9q42aHhdoOcBL+K3+0Oxwoec4jDEsPsF7ITvkiZEkDRcqB7KiDVadYU5gwgwlk7e
OKfp4HpUnqcVa2ve2zRAlKoHbfpTwyQ/6CqOaR3WFqnI3IUii9ooquUZyA/GFsrb
URdyhHFBbnJ9Wvjr3fQ32bYdZz8h2j2XVqjFR3nNdq516XLRmrR2ASQAU3MaGUYV
/cXmMAyC3HQLgjfbP8xHJSXBNr7H8ivxEZil7ahiDKvLWThqIgEAkt0gw/4PE7Jj
dXEqBWHh62Gr+RHYbzr8lRk4lXYBpkKPYrV5vtYHRSwudZJ56SoogWjcsDxX54Fz
iQNehKt7EiRhjR78e3Xfltf9KxnxkmqnDy49cg+9jXQF43FyfTmEXpp04GDpPBwu
Axey/MVod8IwhdRZKUUCmj3K9E9m3EI89Fh9Rh87zzhRwtKLEhFBTxeT3/bKEa1a
YpJ/4I2emAGPPXQSKHEFtO4rT7WOlbYAhqh/dz40JeASisvvRZ7d3JXzCtbYRAnm
Xyu2MFo0jnNKrHujh5o/1j1/SdqSboBL3041Jd0cGdu7f3FuaHD+rtovUEbcpJ7O
DjaROul8wrS9O108yJeczg==
`pragma protect end_protected
