`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
slREphUWM6eY/3XEPhJC1DhZ5g5M39OMqMtFIexdICRSmsYUVrc1tZOd19diZqCh
le3fPVk6x+xhkO575D9lxE+Vu3qZTO76BCfqGXYtQxK9A1yL2JIwTrVv7XdEClyv
kstPEVnFFbMtvp7zZwbvZ7btylYaIGugZJRUpX9WkTthVdhYckJKyFlvAvTuwx6Z
EEuGZTzO0usfpdNZaWvyQWoB4fEfCOfzdTkHXCVpMqoYFfRoECrHxZY6F489X707
Gn87GroqawJp0wcYNskMNHt28EuC9BeeN+PVBFFDY8c3OY5M+7l9DwIE9ZstBi6R
RW5ObuqeSCb+Fi/EopcrOQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2160 )
`pragma protect data_block
63ovg88kH3jwlIsb1r0HxJ4OOVudT4H5s4WOm493nvO3jzkcPwii0QPmVHQxNbSn
UetlqphgtPbURS9t2GCyLWCZx1dRUfug5yivCWDdujfL/v5s/lSIdxDqq34HDBDH
2jQo6V1Of1SHUAzEM7l6tt5IWKhR9LL7v63LkP9NNg35DBz2OLKV9DcKohIvcyL4
8KNqZX5RAUVVYWRe1YlIlYcJ3MOBNRv0S+KxZqhafRugQ6JMh1pYe0Kce1ymdjOj
a03C6l+vSE687qn5AGvuupItIBIHi8ucj1HPPAupiuGs9dmF1w7Sz9xmQxCXkygV
sqIwroV6GLpiBsmKaBMtEnMIKZaOgEgXpRdy/DraW878RDsIlRZ7fHYG0eN3TkYN
rygHAzuXlDen9p49dqgIWaWkzaeSEJMyavGAOHtF4VedlTKDimGpV8R2WmZElRxL
ymT3hE18PVVG7nhcB1J2oo7b+lE3LUnGKyS/GP+pxpOyjjitBzK2BHtLnDL/6Kui
nE31v9sd/F6CL74y+t2GIz/uXS5KecK+NWpVsZM8FKRoO41bNi/kv+5QudcbAEU+
Dj0yyJi1sDpMZ4RxA6Gw+DrYKWUxA2GPGdiWJJ1AXIhk5Lra5wrEKYUbgk2TKJKA
Bw6nVbKXTYV4QvMawqwheUFTTkhYvozZNIt4MinImweioZ7LYHK4GIcxj/nISZzI
Dmz+wqqeBr4WKS4vZV9g4xTvxUvUUkZxuX5Ww7nw4TElME04Yoccil44J1AzTGFo
3RdxxeJX1LCfC4xc6yT+xEm3tCnYi3rYK2+NVBBKvxBOkTgxk7mEe5Dk59wuIBBG
qW/JoJ59qFF1y66KYAEDsOVx5b13mUSJGJC9YemQEZTru8kL4fzkvfv6RXiUNOx9
RulDYyHZ6JAJTzGqJAldSbult82IyAkEUzLMEzskBVInM4StnwisL1sEIlX30p9k
efCOvpP7otZh6eaPHGY+vOvFTCQ4Mf9GheSclrIpZamIU4ovAzMlP9NrKigFw06I
R1rIV2lWH4U7RGFU3hP6GEXn4yNLWonQnbw/FGMEwlmyzUvX6COPgIcdOr1Mxops
BYOQBpOPquJNyQm1jpzZbsuHn7iDnyLZ0XlGI5A9QJ6Pl6sNDoAu89GCk0ji32+L
ym8BJaMKcqbqvJqb6ukWp1kmHvWUg5oxkzB2pdevWLwxNtYPeoJcjCnxhOA49Va1
HfYcT0qk/0lDwz2HaHVxMCPdAp53O9jiM4YDBUcxkEuVt8qBGRKsGbjEwVG0+8DJ
TR/RXlVFl6Whnb0XfouQzRkog2feXxdxIfY2Yxuwe6EzVdYSN5h3KaeLXAi8K+rO
GCRqaNkvQuvTJgNYc8CsRN9uBbj6T97LEv9KfusTLnJJZ2WAGrGk+waddyZRY0Xe
AlJDtflTz9PhuhGL1K0Chh52wvt3J+FRhkWT857Yx6+v0Ezz82lihuhsV2Zc0Dqf
/U4RH/kwMj3665oPhjFQ6A/7u3KXcNn7hq8usfln9sFJzz7ZWXIC5bvKOZxjZSYZ
xzd7yntgddwCUphXvlFu4LL7M5AQuiKPU1g6ZrAl+NazxMTuqatggSPqosXFB09s
29WQxznASncl/f94tysyfdBdPxbuQl8nFjDpncqEvkWjvLMnrNTJ9o8CLI70BFgC
HXpPF9fH4c2m+rXhjd91+nJITGZBJX81HzSMX1wayubaDRMmwobL3WwLJ2NZBklV
4P21ki8/1keIV/rJ+yv0qeWWbGNXQPYnyy/jJw6JPO+CjxqtWHYjTU0JQhv9OWjm
+soN4Uw/nhGyRNpkN7DZomFPOAK+KTM67JpEE7+brh8WXS/yIqKfqC9ngb9Z6HN2
LzQp2d9NCqT/HD2Ltf/amgazAuxZ8Um+bctu3/Zc1zupNctguBz+pSXH+wAdEA8a
n0wEJpmdJmJNG+ONjt2vuHYeoXaLIUkKNBo1P6e7Y3+fFQePHRz+X6jA1OXpCVeD
JSXtM/wVCpNH8UiHzTRPkL6I+sX47D8DDHM2BjXutDYI+L/koFP8gp4dJXJ0UZy+
hb2sKTVgdd1IvGXYK6+CYor9QItVmWppN19TQVSg/c5bY91K6JC1sZJ3+1yvpZuQ
G7p2HVvF2Z7GJwK96w9x6e9kpvdGlTSM4+cZz7szhwt1sUR+qEZnsRLcKX91ujH0
0iXvo+Tc/n11KFtQ4B8pRjp8u1yHHRaHKhVaHvgtKfkzzKIFzDUDN3lJm821jox9
qYnTbJEMClxCljGs8utG6xzdtR2h/SzhSp0eBoTU+DdcVBOUVv5Qfra4VWVLUBno
ItySK1MjX3txtq7++VspUQ09rG6DBsPIJ8LZ4Xszmnwnas+DsxccmnCp6IWm0joQ
gfQQ902oJXw17XHXLgt0H8pUem45zdNAY/dTqAYkvwuuWwxvueniQZQ+PIE0JUxq
51NQ12U5VISTuFPbit++qCSyEMBSq5rybOPllXymp/zQinEWT1JB3j86dMdCF0XK
31scNMzqCZGZDn5LEfQWkDHwpMVxiDBjf8kR5kVe34MB8Gvzqpz2q1kFlFNdypzz
splkgVqRnxUQ7Nn30B8v3gmIPMQ05Bn+pyhUJ7+ipIQcET6GVMeFYmECRNTPolJn
YxDWT2ytQnIzeN9TA0Hg4yB0uLlkPcKv6yKHMsw0e2e9Bin6H+zyTVuVvPPi/PC1
MQI7XSQ8L8Ii6LAyX0OLL5XlTLo9pxG8p/uHyvc7+E2fmmUkjs/3q6vPFCoiKxTt
lud7u1AECevtdNF/8YJfzQJ9rFMrZZDLNvgM5olodXI4aL2Y5yZlTIJT+bj0G+Js
Q7u4fZuU04OMCUtvwrEX2QGGCtn8vbTDDJSemJbfiCYcf04kwVQcN/SHWvh9e22O
`pragma protect end_protected
