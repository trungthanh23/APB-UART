`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RLqFeqtPcZSc1oq1DwLtW6vKvAR2J2DH5CxmGKGkTW+rb/2fl+yNCR0JazBtw4sX
jrHefUHE07xI5tv8FsWu6k2wCSVb19TWw+wPE/yAbQUgckpaiSI/Ym8oUG63jOG9
hI09RT4f3H13uS0zbni95jhlywkN02na9TZJkPk1cjsLW8F6WUGURsedRvWteCfa
JlVS1AGcQsukSTju9lvbujCECqx8H5V8T9kTQSeYPYT6lW4LcqeLxoT/SkmTf56D
RpDFbnZDErDJGMbLiqNNKjTtRg884lzOzyCgHoWhwZDXGYZym3ZyQslTkJIqNkds
WFcyEwFnrZ0DNTGqoA2DOA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2272 )
`pragma protect data_block
UM30hthbQfafuOrACp2HPClOzLrnufsGim83zVaT9RoMvClh9flAqsulb1OGMtFP
ZkZGb759R7EcWqv0e1XO9v27tklKlpqt5Whet7dREO0LHRjKGSj4od6oMcelRYVU
toVTQ9/5CrxkPMAnOZIlPHRBY5tjGlcb/CRuf52ZXDaDTwpmepUDJ6+wGOyvm1ZV
dhL97N9dOeOYyYjiVsp7EpfdvNRSsfvZuphkcSsaW5Hergn/TbVKe7yIMXkS7oTv
yDf16TEBdZliKftc4tEqo6iZPOk8zbXX4gHr+1tlP7yqtpd3PYbujRPHfmDYJPBK
0P6cV3VxkAsEyzOvM4pP08cAyjpNEfQ3TX5LBta/lFaO48t/DXwT8OQ4aYRjy0sT
nEKfazqdxTCNMzx0SU0SJ2jDMCmbBuJoS7DBwhkfzP9zPYaWuNDKs4rHJ7mB0fmE
5FZsjWo6DLV8/d4z7x779J0Jr3900UFY/I0ANIxEzYtC3T1V8ih77XQxS/OdSzto
MXupeJr7P09rwHk9itpqQ2Dzp6KgEdUk7uOL9h3ea7swDBfCIzMhvIo/fAJEFvYn
1OBZY9J6E2i1uljT5cNIuYmq2ndmjxM2ETCfcxsdeecr/ltjzx6K2aLXmH8afJlH
bpahMcK/pNcAHYL/u4rNTlDjgwWW2XSIY2b0z6J+c8ncasoneD12xNWWo0RBPBqf
ennsnZRksJOqMqHu7JancPxU1LVN/luwuCfpLcXwYGc5TC30j356rk9Cd3c9xLTD
X5SgjBGoGeXTBZ2VYJ/sz+YF7wTDmaKwrTbxY3dC/0ddVOrRYXfrHQWlfJr01uaV
+NWIHMYV8ue2tIo+ZAAS3ARZpSHd88oInO7E1Y9H/UTX1Esn4ntKWUlwWZNEZ0on
gavAITycOjZFItot0zbgv4JDqAqY4aLwqjjCEQZ+4yzaMltL2F22vmgX61DMcY4s
lhuK2EAQTolWHojzi+OmCRLZUt7XTd0YLvnCdacMSklnp9HbQAknAD16Mnh2o6Op
7WByFwWiCushzTwNW7OWsA/Da0GQ+4UfehcyoWaPJSG08nAbWX7QQA1O1Gx4IJUX
5A52QSydRj0Gg1QU6YZgD/bGrFrQO2YiThC0Ru8xunFLcC84gDaDIpTAftAzEjQw
xPxNVekyff84C8rKSAMCQcw8zwcJz7nFwcVvXmMmdxLaB3Mk3Wghf4aZWiR0q/vD
5eKFR40iNirV1CRNgtrR7mGPWrLPweRWwBgjU2Wb/PweOlL0ONnB7rWNTkpolSXB
wo5WVg2e1V3WAkIKeYcOO79ERtgNV2MAYs3AvwQLifjzk+O3Z3R2XRqnJWNpX/Dw
WDIOnLkJcoR7jImhp3L3iEkMEGh9L5kzBBxLhpZaEyzBB9l3kNwEGX5KunCTDY63
Uj5FQq+E6+/VSCLROgI/wjCDRuAeA3NHVWl2TJzQ3GjNaqMmcGGrIXQ5mB+CYXpI
OAlzp70BuWKzRrwWhWI35AWWIsuuIkoY5Hm25Bb0l9SbhJFnGHbt8k9WqaVpcewe
baZwmwDuxXZa6W+68YECHyvP2yve84pTF2m/0wSrX59PRrb4OlPYBKp1X2vhTaF4
oj6sWvu8Q2roIo1MMLafdUxCHMaQqJUVZiPakTxTlOsUM2ZhEBLq0hGN2VD0rVxo
/lPw5XQeUVHg0d1rv7ygBOdmi9UhQ8YK+n6gFv2D1wmvgLsk4oLY168dGrWGOioB
Tdm2knNRAu2nmikLyv2H171WyYo87aWclWEIJ/8Os6dQZZkiOfs1b2wLurRa9zre
OcsOGs69FUf5wrM2G6YKYW9dEJX01AWkg5vWaO1+qv0H0Dhi7K4EebGmmM1fO5lh
Jj8XODARJF8iqDaJd45HW4LhoB8F1TMGWOJ+mm12Wo+JKvoY0dqAhK0wOzADZC5Z
Af1oyUL3rylBS8Yn06TUFMmn9QByTRXb1GXk1hbPDgDRUEu8FCtibo39ZAq83Cqs
mKjhEpBJdLxENqmZNAupJ3ehk0EBoI15/0bnvJ/Vo1yohh+yEr4MXrrLKrEIrokA
CaJ8hLGodFbpov6s8/qbGIPK7i/sKjBJeiS4vyyx4ci3fBAUzUW7iMI5nyMIs+zE
8WiIud8BXrSct662WyfsVTzq4baLwybY4eQWJmRely74A+u+dj72bssZaX34kI/j
m7wyCRFQhPI4Ev0VOChNOMAbssX/6JY1pEeDH9BzRaWQaJe8jTdpQt5KTKb88MfY
W7NcSJoBSZ2zwX3PV/8VZytQ3ltjO2Eh/D2Uox0HoiiWi7G06U4uGn5phyOlb+Es
ofb7c0aIUWO+v1bNGTeVmTfiVL4h26XReRAmDULXLluiasUsJWawYYimrbTlOVQA
x47FZxDwpqLLQA6rdaKFlYRFnXSz+0vxZQwG1PBMSPMqmJ8aAGJF0tZ0bePj8fNB
ryMcBRn1k4K+idIlA2RfzqCA//PQXbMchVTMZwM6v1kLM7fMTY+ij7IgZn1rHiqf
kGDIMWm1Q8NMRq13oSEJc3kzn7rarTHNqgyUgaZ691k9II18xdhVbY2aYiWW2XDT
un26uZI8MWOdnjurDc/Kt5Ia17d/d/kWAvaiU9f02ak1iE15Xm7JqZnk2vNeRy9s
LDEbv4rso+pZAY4pN5N1uyFWCtKwWYlK/GWFJ+oJOY+Qt2IdmkfHw0Or/XiVwQoB
kGbup+fg/6WNeR4q/VaelLoWIgGyAQIgtMei8nUFA6ciQVdtKvt6XcyCoEaQtgtg
6xZzQDBTAhKLBj+Rc3TiCHBfRJvz1NOVryWdvcFFI7e5aGff6lOAkNbaJxdKY/0U
2EnoJWXR2Q6O8UP3EGj+fB3zXMv7P3wEqk+aUvQbNsGFmeB6Qc7Y/7xFk6crO978
sW3YwRIGS/WFwb6MV9iLIuKXm1nU/Mc7R3+BYDapUjPVS96pXiWSype2bNcxTo1s
02C2ofPC/YI/mOTcllJ979cCing17KKBqcG2lSaWb4bQsN06Qoxs27iwZbxTBLH3
tTCGYjJ4AaPnv7tbQpFUWQ==
`pragma protect end_protected
