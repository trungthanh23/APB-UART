`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BRvvEOi24JJ1hgD2v9ffPuMmlZmOCpXyojE7BHJUfEVlpeItY48yAmQ9OWptlYzl
yTo1LmSQVQrDXfo1xyO/B9EcPDF6zJ9xbqa2UdfMh6EO0ZQc2pROeWJILiaVcjup
koDJiQbXSVmXRZvsh37swN4jDeo+PhzoPQJZfVJp9uogr1GtZ/Eq/sy45CDKm4Uk
VzxAjfOj5NSbEYLwlOxQX7sRLzvSCK10z9L/bX8/bU5ST1vjViEHGaHNzedoU/vg
1UVT/McEguR+qatA/v+8c9xvC6LfQBDq0kvN3bxocbZOTwYiY9hqR3DF+qGaMVvi
Dzhqa8m57D/DzEL2FyraWw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2128 )
`pragma protect data_block
7w+h8rutEiDLnSZRYmRgxSHgcxuODVyv+K5LY31yTcydAvpDSPqDj303Au3goMzB
g9/jV8bisVZB3VkYTlWSEne3XhswRCeojeuNI4SIL2T8Gb6V4uuBPKwyp8Y5pj9M
Wng1mdBwESz4/lU8z5OPbu0ciVA3O41RNdCFD2qG53rdGoYMvJEd/0lgDP2URUMO
K/YgyhIG/WCh/t7webZk2Dm5NTTcdRaqtqcB5DmyJZB7hgs+vUh9PxIeZxyXBp7h
Yeihn5HLIGzqIUDluRtB02HPDDDBMCxM27ieXAD4wSyFwjnlxe+2LHUmeSDSHFGT
tc25Gc6uelJGPQ4RSM0dsFaRD/P8+5dla3HQIjFveArmHugviA1DWp1y0siXLY2r
bTF7G41IjC56Pf+ZEgnuLjCLkD4/pmlatB3lhMsrpyDaj0G88j3mARp2kUtYUgJI
KvbUGkD9Jxz3Epy6VuDhRy83STlsG+M+ex225kzjRpZcs2Zq/7vDCoqJHIe7kQsc
TKDd+QqDBNV2XRaSYFJo4EmycrLzxTnwXPzWvCP3XFSzy95WetvpPwF8cs5uwZCJ
eHe8CpI6+eTRoY48UM0lGuoWZjPmWDiOEvbR4crEsn96Oo8UnU9u8Fbvhgrny+FW
7+D5LgOZze2OL3iLJ5jQ5Oer0u/KqjaMQ6gghh/bIxKQxovjCJvpSCaFyv73WSvL
q2E+a+wbZHzIWifCVhUjXeEpzoLjh8lEgJ4jdia7zD/IkKscyI/VA2Lb8nutIOiD
OYSxa+K3frdK78o4BskZAKRBat5SmFLntRu5V725wsEXujvF34Z4InKPZBy8witq
xPGgDfR844CeOVzOuDH7HFoKjdFEPyzIAbIupZYEMY8wDXV/EddF0y0kENLwoMnO
lYWGZ7VeSvOov4yplw6W9EQKpjfNURkyBUY8h1XR2rjY3nVbS1iU+7BHP5h/oNUx
UhXdaNCM6i/og9RXpqO+S0LThyRGP0nd1ubvYOOLuccV21uLzNa+rt5l5MwGqBe6
LtTvrkhPOwueH4YneYwTA4tccn03+rx0QX/+HDQzu4QH9R6Je9ygdu+ijG9Gthqq
g4xXXSiDuaC1/Z5lD5rLy9gRV6/zEo+EHu7eOeLj9DR/nmt2NR6tNvVMlimM1Peo
lmj+q36MdHP5dnNFJq/R/KtIj5HzeHFCb5hyVPn+ZGbaec1JRBChmor978FnIUdS
F+j9gVfVFyYR20WnErXI/UTxgRyreC4EgqWjamvddjIgDOAU1o5rMD6jwbvCj+zm
4lzINuhKBOM8Bos6PnOPwKp4R4dz0VaabsWnNDDa1oyVB6r9dNvmsqvTMjiWbWvS
Kyb2vU1ynKST1dowKmwP8gqXUXIAp3/HW/O37QWyOvnZrmObwJkih5CUy6nBmzi8
XCt94NFstgsMNEcfq0a6w/6Ap5d0X3Oq9JMQsZgsY4jhkPbDRNwkFzx0LyTf72rz
MIUMzXjGtaOnPCAtZzm7qmK+4r3nooQhsoEcWNbHCDtiQf6Hi09a/R/W7lQwMQ9g
jzS1CfmiuevA4L9chjyI2ky+mYZMu24Q5oFnH1Jm79WwMANRveZvz31jdDovvfwN
SYgwyYu/JN4TKW14qn2bA3h8vYzsW7U39SgOHenZgE0AxUO0ROyNZRFBOxPR1HFg
8en1be9HeMmmV4RYsbkt30ywNv8NEENHQWuR4eKVAEh69JUZf6zEVA2CJV2Po9Gu
KWZ0wMxQKWaCV3NKi7v3fKf0Ku2RvF7MjORe2TNBhXvA8KZY0yp+/73r5gFwqLl9
Bhg7z2Xc3CQljxXqrF7IR7K8lefTyVEPP9DshpqisO5yaKinhRLIgaR4NR5Z4Glu
kX/Kr7EfQT8kpaVMRryKEpKLv3l1gQjGgpKNVB0uZbrGGuQGEyJ0ZtilvNwgCUkV
XAhciQWpoQJld2blUU0b7IpiQAoCT+heRZwi3/AiM9U7KyyFdGRMhOZZ7Zp9fsyd
ckLzkxRjby3mDuipO4ABySSMr8uAXetdXGJO+7l+8nKs5yPVc6QTCINzJdzl+r8a
gS0BUA7HB6XRi6v4XXK11xtpIk1PqIZuorUTPyNsToDFFZJhgFixyD4KfSmYWi61
Xm2TTJ0TigiwW81opqMQBN4ZSHtq0I1Vph/9QFUffjJh06Wy+UU1jj+F3K2DGUMG
mSE6zGNGVYwcCQaC8LSr6dX6ByGUXaLnR+c/VbhaGC4WJJJ7WKWaja/K+kXgKud/
CprBeZVqXmwMSeEdXDAwNPOhvLKeljrvFnRjDzw7lkRxCtzI2jW7qgAkifO8lLxw
YqMCSC3pIgsrFx5W+H7UrkgURQunXklEM33nFGsmAneTlmGpQejK/M66t1945SpB
zBxanXxEUHdy44L6SDxPCkDWNy86u0cocw3B42wKn9ulUpuM8iqnDg9D3eGgcygK
mSNNnPBhIP3ZFBMSelhLH5kEbXWSmJ5htgh1ZhGzQ9CaUH+vT+c/7MwsB4x1b24S
GuwbBay1gvlcQkAQijjSh3dNtkdWh9Yal7htXqfa4blSy/BacEuha5f+8CovOojf
JZIfiKPaUW42FvuCxld8XdXFQVXWX7duuIAbptG0heAiFu9QFHnpt3hZiYtibgMm
OU9S4awfOsz7PwMKvbGrtYC84dNlS98QR63RH0RHxtTf2IuyTavgd/FNq+u/vaG1
gs20aCSz1Xgq1c50GuSgoTmXt3S4GOF9WiNby8kwPufPlmzeqAYhGe7ryXMi+YQ0
huxdJXovcf4E4KIPUirb4K/F958L9Ud+pxu9D8zjmtvjMM67uohN0klE3I746HGF
qqhuYLuklbPBxuJ9w+fS/w==
`pragma protect end_protected
