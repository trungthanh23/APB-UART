`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GnW7C67eUzyAauTSS2lf0e6azQCM+WXm183svTeyZ7lK3fOP0V+dnp8JvmhFGQQP
3S9tnxCmoKdzyiqEOJtl7Yb5Nw3Ra5nKao5nvMJz2JIUAGQrId2rL8GDtCxJl8I5
0XMwVn3/mKoLuGSq0gOkyFNG75c5ANirEzWYC3QXCyVxPVf99lM4Y/DWd+aWPz6r
wpMWijG4O1WAuxMcWd+DmIixOQTNiCQueTY2bdtIp1yqpjlVUpBs4TQeG1jF7FA/
AywWD45O8O1YKyzraEqDJZWT3ISrC/eab6m530v53lzD//QhxBRNlwZS2hZa290O
I+unhs/r0C6i4jcGhFCbyw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3664 )
`pragma protect data_block
59PALDoFRdpVSa9xT0PLAcUgpGTVlGpaiku6IF6cIX0Nr0rpuYYAaiGS3tdXCehD
jmihoQ8oWikpPdMNjhp5GNKNRBPwq9nk+DFEsfrirY6ANbWd1AZl9pNeMIA6cuEB
WfjsxzOpynOGupdEWdsja1V0B7gj2Jr4n0JXuwQq9EmO3Yb0CpBVXAu3tB8iErny
3v7HC1839Gro8zxx1BLEEOqIq6B/wNC3dlJ636lqzOXtWBTmU6HMtD31K/JCbqyL
4TU20WxFmxv64PDACZnmO3Mgb6CuiQPj94xnw07eflX3ZmE0rHNasahv7u16NlxC
/vGE1YP8LbWLqLr8UhRdj3ILOQwyQ/ybRyJaaeVccZYSw597nJpD//novax443p5
8cLVQaKbwoxqCN9wSySy0UH/PhLgmgSryRUsNPBX5QkzHzdxcmcx0wW5pFvPIOm6
kqpHuv6Kck1fIzfKYy2+xcKPqNcalmB5vlYjC/DWzjV/066j/z40JiHovQrIdf4O
Ien2GJgDVkSQp5wd1N6nucm+S+Rc8cxsttQjnFMcuLutCzLJf998DBAdkORc8BBt
LOKQjQ298ZJDVA2BaR2YHjgIqSulLEkt20IuzQaNbgzao5J3gMNW4kM94PH1alBc
gRuMFoCq8uW0GtHuMzyKXvqvgBZwU+eKZ56C1JsQXL1tmhYzMSc0E9e9qcigY27j
YfOogza6zFCUSQAymTQ64dMLCN5O/ianqF6q2Y1nGqvW7uaErxC2bbqzpie0mpSJ
YwIT8qbLUE7qO3Ec6XQgqFqiKrE1pVitmoC4TCcqPnjB4XYA31DZ/rCmXCcGjM/I
E+E/EuWY9U6Unk85Jjdzb8Dfl1jlEH2p82gsBakuux6COwvo2UCJDf9HfThzHHC5
UMjRdCLwfRuR5Xy822lnHCmXWV6iAUZIF0aTW+zKBo8zmcLuDvIlAca9M3hAIzyt
VDpiU9zzgdV+RA1HSgokKBwLO7rW1XxMQ0g9H87JyGVFw7gWpVV7AO0Y3oHGdUZQ
BD2R2ZA9NuhrwgbJYpXNGEYUO7L5juPPQY9iVIpKf/DSvS+4VBVS9bnoRwU5ofq/
Ktp2oY+BlyEWwSuUPsYNuuX9/YebVuf75hX95AOY5iPglGyEKKwmkIf24UHhqt/B
yFyTkGYgUstiOHk1zdF3n3xXE/QoDYkoDTCypw/y5fu8KAE3ScTBx6CsRkHYU22C
W2v9GRlG73EVSAxYQJ6zNHF2/AlpohCHEr7XM7Wqq1nfsPqlj2/xRIiDJSTzS+8p
/Y70YfBa23StuEhTfzyW9Hpt1DpfcEj/6VXG8Ha5VEppUeDqKepv1Xrt7PBLKkj2
UABuXc9TSbKXXCOUENFxD7fFX6b73I+z52Pn2DmntdFBxvy+pdgAPRqjrBIo7Kdq
WrMSBHq0fA6jyeIQ1UZPUz/l8ijEmFavGTEAgdZiwuSniLr9ZRrCLc6qjfjBddAM
aMsmp/TP57I6QKdiS+7jj/O4LNEJlxWvALwCs2aiP+mkJ3TpUjpCzvnrnF4P8lHK
rR5CGhDmWy1rbnXeOIjqSx+rvCa4wEVzbkQGfFWxN29UhL5KHDG/5VyNkHSc0ItS
F7upu73E6Jffd8bkX7UTCIKYMpa9DT7RJrsZFYzUxBpt7w+GHLsENlP0W85iqaVr
/BrQNA+DZslQrq2GOQ3QQ1I8a+jAS66XU/zK0QUb+dC0WWGLzL80YyhIA2L4Vlwg
2YZQhU9acZtpOWZxPxLc6I95Q+0/+WJXI/NlR+TdKm/LOPwVz/DoHz9g5csJ7ivh
RYRaW6XDaL7t2AIdSBZiaBDEa2cdOeElaXQ6r/DnwjFCJe2zhUZ7Fm7nxmKHSBUC
Xs9ryJzkxOHesIOQbxY9n823CAAYctH6n6pXGva2rgT2YDnxlTOWUmykNHhh3MNm
v/VPYcYCwPiT5VDGvwVwMBN+EWovDaQvAY8q+6aCfdKh0mpmqgaE9hK5s1PD9J18
FSIa47ALrdFbCOWgIgxyGhpZyWaC08jDR+3JIPkHsC1NG4kz3Ry1CM5gI6DStG3z
aaWxV/Lqx2CJ0Z53Dl1guRqam4KcMKVhfUHDNgjDKZk9erq+b+uSZNyzotqJZUc9
9Brz+jXA+tz/tJ4iJ4fLgoXCV+ClTxABgt6Db6cUMjYAO5SOn6tx2iU5ksteCwwf
nkRkk+MAFWYwsZLUaTaO5Ne2xN4bCCCyJvuwMSIe1nUD+edpWZ5bkIavBZrE3Phj
at39C9GYZR6IAFwHiF+wimMjMRi/E0fpoFlCJUz21hXtPjbgayVoezc/1XoRNClB
wVm/WsctQzEiDr65qSQw1FFEfp6zUwwRjpDZ/cQunas10kat0aLFjoWvYUugq2W9
+GGd2TjtRATzKxviEhf2y3FNJ+wdylvirGjDjTJTpgvdv4Xyh4kLVtpIUI+KyfEs
mOixJAqV9g+E7I9cbrgTaeN/sjjBgze06Y4L6lCu+qoVW73ax8bdX6mBvJN7kykJ
n1Iyh9Of/uuNaqV9Q6fNU4H5ZDE7ENRiBvnhqsFElR4xHzwENVeZ0NLWR5RejSVS
PYz9NTzP3tcNpifrJocHAJk5dgLCtB3x4v4vqbFiNE0haBRpoQMjVuIsyi8Ehzqp
E9D1vjNTK08c6UxPtQCEi2xsbZuSErVNgDvooKLAVXH1Vd/CnYby1saYtgD39wlu
Ptotic38+RAP9rYRc5daifnilCtFbEYDooNn4wpuGIfA6FVBoCWVLsuKhXdwV5lX
Ym7DWMI6Wtk/bnvFnK6JZIbHq2HfwpITPyv70B7z/wKfHQqeKivANTAz3hfGSkOO
X3U06KOoTO+hiaPLFJmXGouKDRc/0wrpiL+860UJhVPFV9xQlSNT2j485RJJtPsp
JKs+p6ZDD9USliNa05xtQy1DD1+8dPCXwUwpC1knKkd5sboDZAn+7NtJaopFLg5a
+aprPAdwWY6f/qbGRsHqdaV8IPP2ug3wf5Sy90k/04ldrn6iKGAziZ4tp12USR1K
0SaGAxCoOy5/Vutd3PFaTaFN8R7ngW2mzsstiD9ThjIdn85UElRsFmvSYMPmguwM
3QqyDvJ7S5ipKNcD7CfA2LJlNR8GlgUxk9YkM3DsQXmh8Hb0o9vqQm96gWKxDab1
6jyG1t7Y0zQ+C5uwc4ioRcxEC/ZlMrTB2RpwiQRRm+DqruEKQUW+uj45wgsKB2x/
RWqgC0w2hjS8eDkYsjpix5zu9xKcPFhBlrSwE6e0yc7r5fBpl1w+amsHaQr7JAxe
s6Gxe6zpZQeFkySifr1al3lxC4dK622nV1GXuZCmUD/GyXfNF0jOXGkAHk+RLeYl
5XUlm72gaBiRGQy/k9GfKYa7uCKzGwJmvrD8N6+oQLHvRfwjHwUBgdLoV3/CvUIF
gdQvyqMPfxERNWF1RCF2Oc4L2traA/thqHYcQtOAuvH78pycP6qTIcCadjktMHXx
hlosMgfdHDJjKf7fDqCF9V2yI0Ylb0elTvdWkotl/0EjZbRyLyEXXRxmz/S4D0Hb
pP4N5WzFBtt6i6MUVZKrj3tc+3bTMD0gTdPHkQERYbxhZI8CRIOivL6FsNYLICKw
A+2uHSYkyGf5eD4mgWjEyFuuclWJqkH5Z4vnZiBHGAFvDBjxdOvRZGPmU7r3AfUL
1MjcSoArGjflJNQHsMam+FkT2qPtiN5rUD1vBp+3WoTcZyRb/4C4f4Z79Q2ib560
HIK6y0LoYEcepuhpY3EDwzQ1Q5LMTf99wGxXIkVLjycXFtyw1PUc07yvPyg8jB5R
JtnEeg6kqzCY3APyLiYQcuwgjjmEYOq68KLdb8eoMFdxFcxG6VK8/2uPerwyOn+k
Lxhq05Ty2u7oi6RPzGRQjWveH7Q1cO2kk/4QJRPRlLj9OiiPUX0ZX1LFA6nH7M5D
6tEUa+9bB3Bm0w0nQp4JqTlErr/sT97TTy/tRuSvZebF6NRYCf2NI3MZ4OCyx8dd
DodoWrb62injwHzBf+QualG8ur2yhuKgmyr1/qA23Bp+NDccZiwmE5sQ92a8F/b0
ioOqYuRZPQWx2q0ZkrKc3FrxRBvMJBN3GSSAomnv6lWzKHOvcqrpSW22g/Fn2sVz
zduHqGkbF2po3uwNX1Rj7UoLXPJJAT7MKzjuysEL+FIDGv2mCjHfUuD8E6L8w24/
Y3mIJ/oB8uvB0kr0PlDShb7Vbqu++LLuIN3S/mnhoPsGVjylnhW5CwiCHV/G8K8s
V2P5HXIoLFD+7UY+fm1ZqIoSJgU7rkdlLKBFldO60G9BkMropB/b2DGAFzhxrAtV
lwSNASo9Hdcw0wipeB0pGAc+2sGwI5RCzi4bcU8a8seokLDBvh6/EmAmVxu7X9dN
XbEYb7RHHW8qbzIBo0RT3IRfJOzG9eKjC0reuUA4LrP30353iyzDZMGbhJjVkYvZ
I7S+unYQdhSwhszaGIRMFe470vh/S6sFfZZeHnUooT+NspnB2BndR1SWClqyak2q
NW6Y3IHP9tMbbNS+/rCEFbgbpe7eL59Tcv5kdXZrJqD8wx//eOh1eqEsjUPGmFf/
R63Cm2awWf1Fvw08k6FkhcZbI0fUKDSyNWiiYbKKE/Fjv4cqRA7rT+x2MQyJhuSx
muIBDKOgEhkUmN0I973V6cgR8JfimcexJwI7368meUZNCvzg7RcwDQRC7SN942Sl
yuKxX7ltjeCURbhVA9M1ZPZfkE/H29+6S4/EYxNA92deCEutmCgmKC7g4YnDmb/7
j6IzOUmEQqNdwDcfUN3B6E8fIDE0RGo3B1sdGvRdHpCV1qANx/2uXMEE6HIX6MON
SrbmxEYYl5QSUDlws4JKTx34tC7qJ68mUmDpX3C8nBigen3bKykk9Hstit+vEs/9
kqzxgzUaRTenvB5dvShrjQ==
`pragma protect end_protected
