`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
q9UkE3aHZkCONm5BEP+tS3ynJtO7BeUWcmhhDDE2PbQS0EXOXoTcQg+hpLwqGdEo
cEO/F3TwVEYY5E4mOXq32RY2KIk/nQPyaZN8YItWThW3f5n/fyDjMGyRKwVimVev
csOQnV2VOO9mi8js/pBK6OVmIjoX80skTZ2CmWcJK784l8/Idp6QoRieE+m2XMnh
Z0vfYjeCsNCMWbOL+1KCRUn4GtbWr9s9uR2lVdjB1ovjD2hAvnrzoQqd+W/0DHrC
oZnag8xN8KPu4CmLT5XWjsAVzvG1gA46LTUEckCUXvkU1VqXatEa0nbgx4wqG8p7
1hsqNCDX93JZ0PGrfgDhBQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5520 )
`pragma protect data_block
fF9+nYbNjv8vlVbfyz8Efvh2dmwo+t074nWdELk/3qIv4dieyktq482UxPydJx8T
VUE31Iy3u3DqD8Bsh5k+KqbSyh3jp+EolBP+phtdUuoGAjhC0B74/ZCklCHCtzFI
0dyR1VQpmfXv4JNLSuc+rSIQl2lfKFrW0hWdqz3k9EwWAyFKr9iq8+DCOMS+/5/k
MzQce5Jz9pIjp+RxSHzcrkTle08F0Vq/pKv5yx5cM2A7FUj4C4aaS8C7rQxCJJyx
exzSiTHDPepdbsSLS4BKYVlLvoKxJDwCYUijp3RqCBpOhHAkug004z5RwqWLbMM4
GEsGyyx63ZNO8KdZGqE+BvKQ6mdgiwT6n6aa58YZCPEY+lp75d6VgYmwmBGVk3OG
mpumoCwSRsCKr9yfpE2z5+zVJpV6HsZnzd75FFVAxNc3AD+c1IfOx4rz0athwNBX
I3ZWL3Y5vUE4C6WemDFb08GBz6NOPVwOZQL7rE7T8PMIviOryt6YIneA3BjjzpyN
rbuvcCjkJJe/KCtkrPzT2fk6idCjvQ5d5/pH/lPFRiDTbuGAfs2zkDwboWvOdqPP
bFX9UwN/seoHZk+2zIRCDmnrI7PxKIMz+EIcx/Db+tjgispyj1vk8sMGFwULOkrS
I9M28aoOEQJNkXHoDCuN2CK/H0sNNd1LomlBi/eNYKvXgqX5Eqzr0yF44JbYj+lz
rWmlFI6NDMYJTXmsTaXKAWEzqDzurHNzMK9yYEXeOAIGps9a8Ku3f5vTGRmxQZ0x
of0i99B1UuIs2AHjDz+/ZLGsX1vkhcDRM+EluO9IXEO/sekkV7jC22REdFR7r/W2
vVSIfSe5AQYwaUUPC7/iPNOIHSwvNP/W5PhUFjAle7Ao7KX1vOOISFeobdvZuobA
nBj0Nme8anGDSqdgC5Hx1y3idKrKIIz1cHgE2ruxj5XVAWVEUHuMSD8WgGvCCVmz
YmuwXp+2wBQ81P1FLwWOz/ZGHbMsOlAbJTSMeQCoLM1YiEJapFB7abor/dPYtDpD
2UZcQPM5iG9tkHfKTHTS+PhdMgn2ZUQQMDOW7wErjzE2MTsvIBsbbdlH3YrVtxhj
v3BHIrWoqoNXawjcaMBPFoN2P88XsGbDsN1JsUfN21KmWTQGgiNKOxXFKvBlJzJn
TeXrqUSa0VQDkec/TLwNqHsuXoQL2bfp/+ARwNuhPgrs6etiPNtXsfDIxcqUGsBG
ehDoOqqMG1hpV15EPAAzcjzfICJQtGYkiJNL+PSjd8T+F+RbGCdNtdWJww86BIUd
DDJCVhY9hB6nfFoOv7lI2H5SLOyuiaEG1RH/l0JEWkf3a3oJKAAlyuapDZ2MXaBC
pl9kySEcJHY3udmxdToo8iplKMO7PlvPODdhRE+aNjsXwVXEK9xOODyoUXQXQDn3
Nf3m0nsHMWZWk/pDTDQpT496VEX51xBvXyjJSL3wymQ0g6W4j5XZkxCo2UMPzTVe
gecxLYWQBRAjkmGDJeUcqvz735fhLcsKqToSi5vcikyl9b/SaYpJ1MzFlnrDdGPI
oCH1ZHcxvLra3zJXoPFVw1tTJSx0bTTTUoik9g/lN46A+owucwrSmQ/p+2dbowxN
dY/4ubk8B9bMBToaFE7On7Xx2WnDu9xgcIHIOeV9QAtgJtZK8W5Ahha0Aw829sFR
Un32ZVKfQScyCKOfKF4jLORlfKHMvTLJueEZLZv2ClZnNb5eU7cred49mwoEU1sm
Lc9jjfz3uGXtCqfWefdHWi89m90Npkg6XjNb/cL0K3bUyvGYC2fglqrIbExX+dYX
/5xrO6UKJgikVCarR5i3GtVksg+hhPDBOM7SYEIBSkje87vUA+fu0ihqnVkfpooF
8iai84fUpMyJwm9Mk1paARSAH32n/m1ahQVkuEYFYr5/k0bZjK4md3Thc6d3+KEc
tNcSfMrmtw6xo8tubgNT3KCt+lOY5DzOyyOqjf67WuQEc/TsVkC8ryUnvSok+wtA
IoqkDUczx4yWeNIcV4v0e/yBlTgA04gLwUalhvuJVwjxsyeC93CC7bLIOz6MWrZ/
s/cZRBCrhN05ZiyGge+yjjC7e2+U9GQEk5vYXlQgUhKTd17SmBz2nWva+SBWZxCR
Stkm9/CGlJXO+ovR1V47JGt8kQX7c+FEqBjrohRBSqi3hFBbzuiIiJvROjP2xov9
slqm2mrobhEcFF9T7qsobxNz0PrHM6FNlic/J78pgnrv2no7ulRDask3JuuQl9iz
0n74MzFd1/naNv1oV3P2aTGBSA1k80r9GoS7W9dZjJZ2BCyLlU9zYSRjHoP0HcWR
eJv/BF2DfCDo4Z3yYVia25mz0RMp/j5CF27skYZYTS0jLiE/WsTCsKQ7cF/JVFaI
Z6hBhiK0IUA3IwOJBPF9Kmb2BBkDQIaSRlVRk7XAoCIwgdnyaj46oKrWjZVO4iBr
nhHmlZJWWnLswIyRofR5m+ax2BbZ3x91CHv8WghuIiWj41dTMtoxEIocQMO9IL57
eqUSnCyJJZnkZLdQ2PbhaYkz+eqxqHCtEE0xX4myGu6+xdNC2btKNtnVf3mCr/pO
7kncADbJQysh960JKZjrJU7qRTiCiCA3pxIuRXcL3Fju4mOgq98xXR27p8T3Dcx/
hSyquD9YxGbhCHOtuDG9ya1a9TPItgz7Vi1HKjoNjIF/lgdIl+zKyGT/s+QQOSEc
JT9HHcMNvCRO5hVmw6Nq7ju38MSdTnzfE3hXV/39E5AUd1R0SiyR3QRdWQ5DyrtK
Vo6LWAyH9Pfgd3iVifJJ+ledImTsbzyl5opad2nTfujkVlg5XQyLaXyqjLFFPeFP
EFAurkMplNS6kQXwqZupZ3hFlWUWL3mmUfNzbmDQKaP7jvmuG00IcHfbWtsdzkI8
c/ck+nTypD9TFesLHAGYLiZ3KwojZC2qGAcU/8qxqhi6WnzFfhePsTdhEiP+59bm
Y9+jj2Fv1LYfyYqXlv1bFwGjnjLlF5BRYqg+Q03OPOjWExBlnJgjRa1zaWsNGlQ2
A5HLxu3wQW1ymezLIbMmqDh/oBV+c2xlOotaEqJn++Db4Ou44QIHK/Lmq5dDDKeF
lG3vwlp/ulpybEswCH5yhv5AdOf86tssO0axWhkk9NwEXSW1eLceXP0Yb8FN+qKF
NjX4kSWEbigUwYoyPUNIxnjO5XZDMashcFvuifPg11oLjnvvYhF2LMAsUZlI3hyO
7rO4jFgZ1HKYHHFGNGLTxu9t14GvKvJ75LeXXa9Cx13+ce6cRuVrEihVt2H9+jd6
XwuurZUmVzTBPeRy795Z1S/fQEhIwBUsgcIv5DOxsrl4sbjmMpXtWGrDGLnRXSb4
2/Pxz3LiBbtbslD+21ecloqfpUBEGA8fK3FYvlpIgp9HMyRgL0csrlB7lBi5iaeQ
XD0daro9Y1ynUUDwa/x6R+PZs1P83BKaHE74jDXTLMrI8J3YqyugiCyGZxmwmR6r
8hT37ovv0tm8gSHv1UFfIwZVdyUhUN/XdATi8bpoY3aFWmxjrNOYoqPUj9pkVyix
maGzOp1oQhGJsd8krFG52ZEZy/OlhB+Kfeo5MuLaBMBl40wl2tpzRvBB4bYogq/7
cFHOy8OYCASVScOdsOQWX42U20m+2ibHVgzn17nP6poYfc0DyrPjVWTLc8kEVlzp
vqxZaxWejqNVmrXYj/nffzLivmr33lJblIEs3cBTY+SXNkxjuiEPCakkHz3xjkXy
aW8MdbLlUY9nuZJWeqh6zgA2uV4hUSmyCFSBFZR+AWiX84f2vBA1kj2DYbxBb6bF
LkSIfh2YnvfIiGiy1ouHsl7fr3dUDGGg+tJb/OldNijHwI5edJBjDsPdi07DmC+v
amoXsxx8VCexiaqvvki4t4gZlru7ooaiToxv+CCdSzo75Py9eWem0y0xojtBMVVy
jMyNlVDDh2Q1WNf+NIsS5O5mde0eCTq2Wiw5bScCkCGRroaFw2RbN/t6k4WtecN3
STZpLhQBto6vpRo6TjlqDXsS76vKCgEOpIm5PvaKtmuOXZ9ir0Ja3p+2PYELO5sc
5FV5x1mJ6H0y6QqU0+2bS2ubVi/qLZDPWIlsHOdqDqEV3OuxIet3lWgC+RLjOjat
d4QkazAYjw0zANan38Eg/RneYnfkNRz+5mkhL/Wi6UN14rH/vM7hGRHkUiI6m3dk
yIyfr1c51v8xw3qUBQohfVew4hg2nFzydjjL/1att+oZ+NOJkaShh2MjH5SVLHiS
j/tOPknR0T1eOMPAPxE8CrH9pkxzg2UDaUuCcG9EDISgHImiofRCcmBQQCMb2/4n
rAmM1yb5+Mzdg7s/JHzBk3evpvWTNxZ0lOWjXL+xkj4LO+306XjnhLL/6oCNQRUv
AJcO/NLOAny7/7hJej/4HYT317ecX8/XUzI26BDNs0QJsk+8ItDn6hzrbOrCq1pa
WVjPvls36tpPVoNz4ZhMYg/IlDjOQZTpddFSz/ZjsVKiBY1ZOA+NmUsHjg2Ag2m2
/X4+U0EPmKf7DkoJ9gjZDQ22Xv8Zr+X7Gi9MN5CEvFOp+U2e5E3k/8MblaC6ajT/
NkaJVMMLP10Hvz5i6pWiea/DaG1UP6fYjuHCEpCAeGM3yAdiy5ZUAkNzdyk0hw1n
/JChEvsbMO2JcU5bmmDChRuASUdfRCJYtVu1NvfMInCeHMBLhsitXaIG3qw1B0pz
iE+KI1fKNmSFmnSsMBQsz9h8zRLcfGt+DwwpCPA6GGqu2zpP9EFa2pkbbPdSElUv
+yfcYpG0cPCmMK75Fk089z5HuBe7v9JuMzBML7TxV0yzXtu+wDM4kBlZ9zzIRR09
rF7N4iC+ShGozqLFzonc5uFk5ZiEpdWg3T1K36dVOGsqy9wO7Ank0W/798OkIiWQ
jzEsL3SkIpFzYDmkXN5qwagoECH9y+XJfK9wlQ+MK0OqmXaxoNr8/uYzJtEleJ8Y
chM49h9SdGrcK+YXkQD9UwZvOioZXTJm5j9Gm5cECSQQyU/36ghZqDVCBD9osZ9U
GAjzWdsfNcDeaV+DoJKZadEAqIfaayN9Fd0ws/QRMwQd/MAdKDh75o7pONbYVix/
Eo2kd6SUD+S7aiFDo5JbcDOBhNwgza5h/rYNxtdDd1gXL+zx0y9DRc9Za0+kxa5H
u9nf0FYcKF8yZdSSmxWT1Uy+Z2hZOiq0RYhf6AhtiYLFD5KWkv3+ZpcCHxdypdtO
EJOv/+03hMu1vUsStqHSMNF6Ed0h+rsoJBGDHR2ho1mKyjOzVlm2uX6LZqnCo6T6
SdfFc0xm18mJUHp5FT7X3a1G0amH/NWUg4FHVAqftWfLkRSPvAqJoB2QaPnhxi7/
iQv1cEYSoJVyHEevqG0bRExBmOzBqWDHISb6cDP+gdHKHzocS2e9W/Wx/Pkfl6US
QSv5CArq9k4eCj5eQyWYGaUFNmOdjDgAHnFAyl0jC7ptnUYtLIowIIcC+mmeOdiB
0nWbipoOvcoOIYFh0g94qbAQBKKs6T5FzKZ4onw8ffdjjJ7ppgZhtLtU/iVRlX2I
h7vXvEds1wvP8Hg+GjGdxkhhKMOsSognycNwH8G3pEFgM/Vc3yS9tqTlaFhUJHFx
yBHv2jKDxhkEGn9hhg3vS7j1kITZCGfrsKIw8+OFQ53APGvC00+VnCJdMfuFMHLt
elPI72fF8bDDuXZTwaGB6msygWoy2yloXF45/Fs8JQ3+Pe+sio98DKuMiBJP8pzz
y3MEp9mMaLbyyoPpctcqJFHb/XLOGw4y0eEIe2Sq7jFULGmkFTzouC85rv4D5UiH
2ScV+SevcxF3RFB/3SC1v+SjSsjVp51W0kH/3ZFblIL+4XiL49WI9pVLtKMHxkJ8
TK1I6DchQzkhee9SYrE/H6rQT+mYrfVsH+jMuM8wAHsnjFlt0311HweLDhvmfvXO
giBucC3Bqz1rY74uDUJ1G8sRKVBrVQ4R+tKs2Ol2g/SkEpHv/DP9cPkj76pzzc15
uJgRlOUYXJuq4T+B6CF7iYXs/9OnFuom3fQmqyDE1lDpJo9WjAK6NSC+br88lOmf
9f3E+tknScbzmrDvqQ59G/l6MUv3NqUp5CgjMI3jELKbeCLi8yq/7tT/AykicDnN
BVrcmlsyMv1D0FC0/eKZ7ppGzlVO6oZdsRw436Q2C2fam+uY1IzjZZgPeAU0Xh7C
v1IfGeIBLzHKDxLcKDPQOc4lKkrd9zhEAQa21bF5rVn926dmYcmMjTRB6XzMKaQ/
DxaeTMU6EeqO4zXpSO9hDHlOZANRidJQ7r1IsfAWpisVbQudzq5bhcQoxJDP4+2T
Vu5sFhKhQ0dkLgKGI01JNSIZLIuxfiJYW2UENPMLL6Bqwgz66BWp2j3D1850RhvI
/1HM+QIXmbU6NbucZpICaO01oBoyQlqJG5kGKg+DQ9kbYT792chYUOXZXmaVBryU
gubxrLdaQ4qMSY6UGma5czLszojmckhlWGYdU5kElL2MkSOhYzT6qP4LNv0fT1G9
sAzvBZdxRYrcAtRfX+BQgIwH7ntzRRzyhSopJeGXLzb8JmK8LHmTFPmDt1rVMCbq
LYY+1TtC4iM5HGdxgXX5YINlKlcg9G/khqF5tz2mHMU69JTIWIrxAIyi2URW3PNW
Q6lTQ+hgNGQlhqT8JX7etlsNdlGxGGsq3LFdpc2/YrO5zRuBNJZl2e1rqh4tzCe8
ag0Asd3a5FNWQ3mmtCwSwgibSniOVvH590mDwj0Syae1yn8n+71lzuALKoz9v9UM
fOleY5oXHtITWVPPUdw+I396dsZm+AInmq4u9+KEfLYcoqgXweyBUh8XjwlvtZeY
FrqlKaJwaqkLgPVpFdXrEHyaG+rhz1h3JS89B2PbUftZFLzrv9fpq3g6kn5zJLRG
HPPg0fUSD6qvd0mY/IVB47mTyRUAk+/zArc2wRSFl0bmQlzFwqrTYPwbSVK32C+4
iNrOeCN5UwYxhEh7X9Fru+MwABetN59g87VaI7Xc9VnH0kFcg+G6j2ZM/SHUgtk4
yvJ4uERRnPolvUustRDIF8hUI/0diPLkJv8T3FIOHzxFjc3HV/LOh2gw4/1SPg4A
2KyXfYwgvx4Pda7z7TddvB7HBtdPShwwNQOjiYbmohcK4R1F7CltclE094cqL+Dc
NfY6+q9+DaPXsTk0NmzF7OutYsQcxuKUIWf3AfJII1XxSzd4kP2QwWiM0ThW5LWf
MFTCxbvIM8Lkb57yomuG51qjq0sWh0t6tlNrsL+zWDSpxukFgXnktwqSKu+ATeYg
HyOlRuCz9rxye5xTS0MtfnNh7gn3oUS9XvXHVIlYvtQ0wvgRc+D3i85d8p7OMsx4
3P/vma0pnOPAVGCoav0o8aM/X9d8yYMpzzW0t0ZHUghnFplK+B9M8z5n/eMPV5uJ
`pragma protect end_protected
