`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
oDRpAnD/y8R9Ue4JdYt9rs9wOE9z5S+TONOuyBDrb7RQe/+vS0UOEtpIIn1B113O
BxjLYf+8Gh/myqt+HlsZHklHrXGSzBa/QYsn/VfwMd7DA5YgV93p1dvHfoKr+Qox
jbqgeeEopfFG7xbdnMmG8MC+kpUrn9CNg8Psn3+pEMlZ1dpr1CRmt6hWWdXe6VYa
jaF7a1yqXTjwQMBL4K42MjHaSlPSAJdV1quXCvaFKBVb8heZZJAfP9YB/WcCwLnn
X9aKnTwxGlZo9H4i9sHSC8p5gzx4yWbNzbkIWIPieZgk3VVwx4OpzYjzw3NqXxSx
NwN+qpo1M+KAJJXQb+Z1RA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2352 )
`pragma protect data_block
SZHQUFlMDMj3HQlr9wWIEjM6LMAy0PKVANO3WP3AMW0uafi4T/cx8p7VohbPPtmM
VRK7pr+by/fYqaPyl0Yf5iNxsCuSxGKmC+0WSCntUP9+FnjQR4rY7pvke6e8pR/+
sD1JJkph2/97a8QEPCj0x+r5vIPYwLsKLo59+FGD+TYrH8DWfknMfz71z50JiaHF
rST0NfPGlI45Y+3ZSs8cQwydXJJZcBVuQodVFfLTW7uAHAoIlYr6LqDrFiMafpvI
tfhAiGWrMaZ6K4aXBsVDzs7hmHJbrN0O7p1VyXPPdzwX4O3EQH0q12JLS8BpKmwf
dVUTZppKsjNFliWuhjqNqznulEf1vctbx+toFDhFPIRS+ofLVzIDgimD+9W46CLB
X1xRoqQiOXX517j/V6ozauzTatDuXXGsZtEojb7mG597+C1o1sz8lDKmLa936bi2
Hsjlhi/8nEGL4IX/1B4LbaVz0TYFYr/JdvjEciwxBLTkuGLIfyuvsUixwSEXW3fu
XHOcGCp3uYgmRVPhuA5ZIHHaOqgvAQjoit1YPeEowUe5q8iUjQlbQyYai6CTq+kM
RxpHIbz9rVHVWbkmmObArNXMQgyltNGUy98M0dRczoxuDHRpbhgrsBY2ur5fXmRk
+QALc7JfAnuNG2SjKt8Oe28515VSylTGAF9K7HUcX7VIPSKW60ttxzUMAVzacmqH
kUwMRyxDJswWdZTl5i6jsoZrRcunehpZZ1a+G8wxv7PJk+9AfUivKrtJN3Dk7lhX
oND4Qs/pJ6dFpM6tcOPxzviLZxcIXc/sdPoNvCHME15rCC0Gaicjys9XlqzvoA1N
kz9xqE80a1sO5zOepvMuOfuMA5wRvnq6Lkrr8VAMU8IW0aOaA8NZjBGsikMSwjNm
lK1rGGUqKCaDpm7mIBboaeKYXi3jggQ9Z+QfsgZ5B1fY4sJwjxtHjN04AK2by9je
+LhbaGBg9ggdQUBScsi6iuhFAf3AXRQ+r3N9yQYBUzsxg9gC9UzuTAhu7oxOUIXe
yujbI8TICLoM0JepUFm5IoSu5XAeJnKMqAp3F6FrCOl+UsteApZyZ9xVL9olzcC9
8NDi8RYj3cLW/Ub2/uuEmduZu02/OKnG4V9lXF28yqEOvjCIgQdBwpml6qDGdp1T
6F1b3pal5HZX2AVN3nG682F4g7+mnf90AQ1iEyDvDwOgValuuMT6ug4aZr2Q1Uoj
ACDVtnQa9lT6tEJaYQpBjaX662a234lDQUkomy6kl9kjDFhD3B9GcRHNIac8yS8N
5RYdMJVGkqTjK78///riKS6dveYzNRNVcCLnHb+gTdM7kHv1BbiKH5shhFzJqeX0
JGAmUfYYY8z5Y3CKyPP/oS3rMFA3bLhYZeLqWAEDXcnHicdJDZ/ZVb54BT0VJPJz
WNKiD0gPIVWkmvt5GVTqkLc1yB8J+8mNCk6wEVhkccRlGmhlmU8yH0cdeXHNbXoO
u816/MjewHnEBF8JU2c5QkmZZmh+GBNNxlOq6gkOMPfqIylOP24yODa3A4DOPNld
yh1fmPYxSK5pDakXIxQ2no27Vt0z3sHdc5QmaWQR4eEIUPYXfkVj6O3aBDqg5S5a
3mOLz7ObNCxtbnoCzAw5TBZtm1iipyFKHZWddwntUWyeu79ToiwgMoqH7qtA9+JA
IVGCc09QdTTk/Co6vSZOi7Wpju7AJiKvkkFoqd73ayUhBi+Fr8pBTcxVKMhd68cE
ffWqCTzjhClSKUdMJYQj6oUKfJJmiVhZ3IIM0roGPTNxo279MZ2UgAtnGiHXv0Ik
D5WBOiS4By3IXMzdlMbQm+GKxvtHy4njDu3oGgoLKfteCfKPKnMkYwo9YLHxjiZR
UYhxnwKS+49b+HBWXV/zNPo1GyMEaD+4vO+9dCqsQHheO8WpgEay2nDmxQa1saz8
vL7w5gCgkh2eBIGZFzZerhFR0jke72cSmwngNd3trD45uRyt/JGh2tfaztBK9rf3
NQR8fAptJwY50QlBydUJMHO7VccWz1N21em825diM6yKQHQif/05tlSSOf9sUaDW
AlF8b0Ht48QJaUXDqoQZeJsrzf8MO2ifn369ef/NR2fvjDOpmYr3MmpOviV6EtdT
L4lU95fPYHVHXx9KxokxrW78mIuGsyO7rKMoy6y2kUN258aHZQK5o8V1g13zvZ+4
nEQOlVQQiibzsA/aJMKwdTcht9/+AohsMcAyG71Bupua03OcwtANNSVA35XnWAYf
oUNSBje56wbNLSLdaDkiNPG2m2EDb3fDbT8+70QWY6wD3df2SZZ6K6KMJLL2hbKl
mtWUemECRAxX0Gn66plcdy+qdBHBx7o0FmGcQ5VWaN8GxfVjFx04AmJpZ/ciTpGs
kEFK7w5qZ00cduwx0/X4F8lkgEKFp3FM+FK5BfEWB8bs1aRs6gjb5YuMmhXywQQg
/I5mUbSW+UkmDxo7s+BdylpwQ/0oP8Z4tzhxA5+iHnVCYQEX4zN6t/dtF5O/7r96
kJOh3ej6e1bmcW/o8CalHceH/ZV0j3xBEhz/UwzXIMaXPW0g15QFsDmaCi0IX8yn
6RRPiwkPCtEezMda3AtlUBCnpfh0vRG34eWOe3+oCngyGaE6/lPOTBubGo/IwHQD
nyea5pdkjxhiizdT4Ov0qjrjYchPAzJ03giv6Lte0BKg3fdbR61z1C7wHugFoRSc
qLHwBSXZ6sI+oLQ9t1h7Q+KjNHxaHT7fKObCnmSYBdiQb3ip57CX+QTgjHc+h2Xw
VZ0YR3rDROOo4ePXTmwAK+0wex8jVzfx121IOPpPx4l7FNOZzHC/xYLGWllKS8kF
6kH6DO6ZtmlJs7qsV1jURNZpdX4wZuRWGyExRMRMbPScF2JEnJTE2hN7KAHbawyz
4zvmv7vtQO9kZgex12Upui97291CXlpW9FKA75ykq9EprfwYlkZJwN6u8suBn8JZ
wM9IpgkLfYZct/qZP/blLvYsRveYzMTEFgru2qKzJ5FkIhMTivMdcOXjogxaSra5
s6DMnZJrFqlEbmSJlKj2SHGSOUhYNRNL0QeJzRZy26cqbnBFk0lxPvWbmdl/3MKe
5awDcas/SAeLjSD/j09xfvUxABebz9EDcFEYoOkG/oUnCzXzm82kbLWHQg8zuteZ
`pragma protect end_protected
