`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Ly2g4D9NpK2N/IHxOkn49+xBU31Vz7CX1lQvk7326MyZpMJNagF0pofHj54weQdE
gpWdQFHOLn/xYlrlnxccqKOgddQht7inDYY6EmgX337xHHxt8+FamYXGdfb9pCHb
8d2c3WHR3FR67fgusbJjwXB73fQ+cXSCsXJTbhXMtJ4dotByBxFIvMRpGPCDZ7Da
vwvz38MfwU5aB65HDlCYQy3c/PerfahLWJap2uB7HlwoSxg86ypANBwxvKHZM2zu
HPlhS3w5wPOW7J7Ve43lhb3Cf6Ap6hGLjJZTgDPYGAW1eYUuCqdy/QazVUrz0FEJ
7kdYpzxKW/7Iya3rt4X9vg==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2160 )
`pragma protect data_block
1IsnOz71u6fKTzXvb98wgjkYo44jH2Y1T7SAu9k3jIYDxmdsaL2h43CEaAuEugR6
2UICOEASWVAr7YtQakwF021hjN089rAzsnyo+cCxlth2rV4rJVvfvhExeWANRBq7
ZH4Qm+hqPZHM53ldeLWS8SDN6Kr0K/Fps+FtzvBPqB7jvChbAOVjF9+Jjza1mkxs
3nkjTPmu99e5VLi8DFwUWFIpSZlGGBHfMyTftxw7wyD5KVH6BBthewk5+A2SUm85
fuezV2lC7LAa1GAoG2t6Sxt4ivc0VrcS8PEywPt/DoMhNPipeeOQVYfMyXpMjf3c
vv79PVqHgP1vcV7yOI//PYz+G2c1AtIq6AANy5y3l5bEBhaW8oTqSe1M7LhmG0yO
3e9UOOJDe3fmwlq+dLuHygF/3znL2wfcUIZMniYKwISsWxaPyzMuAPV+0BH4Ps63
DdVR/F6/OyI3uuJcxVJeekqd4wrrcl/JMtAndXGQAeqKjWiIRXu4TvhoXZnnwym3
oF2pma+6kUCk1cAw5aMnsxSfjdEukc8uixbjQ36cuDLjN9cRSAmE102QERVwK+q6
nTR7yjPtEtOxfGj0tqdEM10CmesB4g76xhWi1CZbO+VkkSopT3Jg1UYc/2Su9YAf
dV+RZEk1ycfd7bcJUC+hMWTxmeec5ABnQ3FaMXffFznObw840jjh5qbOK2VvUJCu
Y9RjqM9w6rYe7I8I/u1MIaiGn0RvUqUj/9B8DCHBN7gv4+0fi541x9l+++9xQz09
pWOcqzzuMoH8lMpRobzUzUVxslLAZIl2znNZzzj6W5TB/ikfZ+hYBOT/5TxrWOmm
5mThGDkS6J7qbSLBUbMmIH12PsU0miFOI/kM3TAfmMuxQGaDXbIohJ4STo6EbLrq
aSCHHJ+eBULNhmzv9ToL9xr+yQefHQZMt0+CkK8jhHr+7LQP7xCSdLpKe2vISNoI
Km5gFWQcJUoMqcKwhvI4BtAC8iB2beUnJ2pPyZ/xlF+UVdv7dcQx6FbeCAhccgbv
Bh1rtBdpqy6ZN6XQmwN+cKZolBegq/NhVaRNMSoTIsrzo+nWY10CtfzX02RLssQI
UzCPKXVPLa1sxd2VCTAlY3yNrWVC/WaPpnM7bbGaFwLFXyHbK4wvwbc0wTsn/bUD
kaqi0TTugQRjSAUc8j9xhqFdZD+ZmI5g7jvgZeaJbjk2PiZBBb2OPnFxxGNBYEIp
ljbZXMDxhH0OI0bOMnZE5/skm5Lz5ZqWSHYHHAmX+swghKGgy9OAHvSErFQjgnG0
RyVIIiZJcOC2IM+A92aACYB/Zth1jxGLsnMGq/KStWQ78OKx88/GRQhXQzhkefd6
lDW4cndQV/bVWKVAIRHEBT0DNTU81cfXvKRhJ16nVpEX9vcn8FGEXjsZSmmJvRtZ
qNMBgAHNyNRvGb8JjnW0yBceeqlG88OOTIHPsp0MSjLHoQ+9eAoshVoozh+nNjtJ
huUIhhruB67SJgqf9gQSO8obxu9eHn7B9L1ARu2KTi0fY6MM4RmRZdwhpaeB/C7Y
AaCnhkLYFu5GeXtrWbD8Lb77islezUN9rE9VvL+ocJb4PiPg3Z0RzczLRuFWIm9+
18vZSw+bJ9BkkDkop5C8Z72dqw0b/rx8Pu81KNJhzpta28iP/WHNjTATF1S2fugV
LhovlGBfQO5kXfinflRaK7GsRaVIWUg3bP/2T1UyV+msyiz/P7+rS1EajVRd2dSm
g+ooMiMLNfhOiR+p9wrOcnKn6Uo0lJQsQx/CyS3JSWZ/lFRfDqQ4b+CNgEzHuKtU
4gd+StMd3QzFeuUrWDRyqib+jRz8sakT0+35gGviN6Iyy00OF6WK2k7f3TtdBr9L
D+sNz7n8QQPU/+uKUjWqjRIxWNRxMR01smYdLUg823I/il8nyFdqkhyLMFK/892i
6b8ke0RM34Xn4cPNJMABvkKKF6PHd0Sk7LOsMdg1lFhl424IzUgLMH8laDAz6qOj
SEu83aUdnzgSs13z2z0P+wW13Zq98b+wLRvD01PAffI9dBAuSPtS75hKDXtJrhqa
RMkeNd58zMV0kTQUA1tw9gGUaeUpYzuI3/mKdoBjqpBWvFFZOqOkbMFRsPu7zGX3
sWWTCkXR6qz8lukc72sHRJnOEcCiZILehqENxSNfJFhV5m366U4FynTj7SxWKY1n
s3ei+xMX1R/27Pjr0NGaUF9tTR5e2HORXEARXU70XqCVa5A8NpywQeKfOGx5eccn
ejWNufkglX+QU2sMvB+45fAFl8iJSnNKSaO4zhMw3Z8oe8wmgJIFHtfW34QEQirk
d3kURg8tqX0RggCTHvJ5cIy4OIedTCO/V5hmpyb4cgzKeoD2wzHRHPu1x1NhKgg7
fqO9W/DEkEtzgRfX+t2D2weadSNW4NtpPZrUN+MbZWa8dJZ3BtpyTocGC6Wu0cc2
MnSrNSOpPuNrm9md/gLQkoUWxuaIg31qAE8A9sZVT7KRBv3k32Ia1xkKccltvLH1
QXA4AbCsHvSJMmG8rOTCUGatyXfknzVy+y7ztl6+KziaK/htF5SrL4l1EcG4fp7D
XemNq+3HEg8UIuKQNfufgzQ/PZdqBh6D9Z7l2UD7Am791yZrnLKw2kaUv2pgsSiN
2m5z/HIasp0wnMr8+eArPawhgLHSIIQ3Hg8E3IscMQ7U8pDa77ucXHQUgt/M5HSS
TeQz1mNF3MBa21z4/wcN0lq8OE64xshcc4/tSlmlbW8k3gS/yJ05j+itw2RKoCMY
sJqvgJWGy0ovQkfahZEsDLq2NPN4wKf0d5RywkGw5DGUP+pi/JI1Mb6Apvasi9u/
6pUSpCCRX8JIh8VuD5mqu83/ZVnJfNFU1Y4QuKjJDaP99PU2V1lyM8UT4etSBePl
`pragma protect end_protected
