`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
n9ITsXsjhDX8PB+Q+8BbCYNfTYXH1jjxkvIPjXV+iHvkehYbdHTFilXUtMFeeT6q
c1gk3yc/nZ5zI4zQ1L4SRVANp7XfePBxGA0ZMtS66gco6Pe10xhbuOMfduLLu5pY
KxWwyALyzykvgYZMaoVHu3QaB5UTKFIZZKi1QX1zpsZ8142sGhNcaIBe2C/XvwtJ
HT4CIUgMiPAMALeq5sTv+W6Z/IYGTwhcV0/b/4R0iDoGolE7jdcCZTBISlDXOLYg
dIVGbP7L8f5xbyT/syUR0H4hFU422qyp8Q/r/G+T9dzyYBq+/ZCEt+uZ1meb/XD+
uC8p89fZTmNAyJL0o4YhwQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1280 )
`pragma protect data_block
BVsMYkCb6buNYofZSVTtnXY/w/HID0Oj19xznKuSmfogaZt+ABKcnk/vIyydCCJj
nizUQX503bUDupIdAScLX07k/M8oBoCR57kMa8H5tmLJt5U7jgMWZXmL52NfMp6l
ujFWnEWE4/0OjEO0Rt8dYwsWwRASDt/cODDKJC+knL/r82ei+21rLxqKbYz9acHz
dsxY9pdrYNJfoLnhlR3eR44TAc1LZCNx/jYoO6EvnVi026W/odNnnnge4HD+WAiG
DVHejM9RpEvoyttJFbfjkSbbuGZ7/7fiFvx4ptOPXcY9ueb2d0dyBainCDnbiXnR
n5PY6KZMAW9qGuyBLQ46rrGb0Iq2sMLrJQUrTzMEYx6exEq/PfdnewAkthFpKh4m
wK7zoAzN4q79zNaxlZURB26cAoGjOTI+FBlb3EAEyN9oIRTx0vx5EV1D0x7EXVpV
KnxwgF2eYWEzmgione5Y6Gtv4U66+J9GOl8QNivSwKS4zri7dYc3LVGok681b7NR
tvqotmbX7mmgjFbrVnuJOrpIhsGzSKNLPLRSQhbbg8b5dDRet98wPGZT0BZxBLzS
dkCf1PrZiDkrRkFVQvi24Po5MoxPYuZOHXm7lAqub9WrKuoa9WPoZN8aoY/CjOqV
0RfNkvYG8AEQ1hN3R5fn7VlK7Q7y8WQL1wrixYQraOtuLFWlagAwYeFUH1GdqDkf
T/MWiWwcMtDIRw9IhCLrggSCmwzkN1tmiSTFInSj8ZlXHsPdXG6ZSIyDs7XsgzKR
0el4WFejHn6oNX5Bdhb5rvSpTmOS8QphWiCpguqVkwScl3kREAj+Ok2iBWWktcni
0+Crr6cRwvsmzvLUl0V2+16iDUjX1RVolkzx2lkVG+D83gZPEfP7dhrNYuQfjXDm
bumF0Ki+zimwEKk1xOswYi62dlVP5gFI5eKUjAiZnUO4lvAD4gnhcaTR+L2VgWnB
4h7n7VDeoQi362Gtiyc6VSl46YH+XadAXQ5Ks8b8VFNJg31F1OM/my1645X3tlYe
798SbDAFJXTs/PtypIYIxTXiYKEYvTO7xhU2LLFPA5eYXlhxkuoVpj9KsYSLIR6W
E9T6HU6L1ggxpyvKDk9qYs6EOdMtKICnElbShySQ1UiWJ9q+A27eNdUpE8TIqvWv
/ggjKGWn4oqfdA2dVJASEApB04Ru6FdmnTtz8Y9TGs6zIIDlTLXkAf6MDTWAMSY3
+GTb70XPtpcTG132EYPungxhJ9QqUbGY7Py6IJJlhX0xDyhTZWrqtmkrOF2/YNKy
dJTi4NfcWf5vOK3HGQ9k8Nq06RNnQ4aHvR+eBpnnLRzqCtC1sDW/PA3Aa6Nh0GET
lDQA9wU/Gw2i7pqM8jFeEyUwuVojbMmJ4cLQyR5TpNqyXYREwYBUYaOG6XGq5O4W
Aa8Jikutiwyq+cTZRzCcEaSdqHBXO0xk3MdwWPaEmCWksWL330OGEgGyiD/4G0ax
NsaXytC4IjByAgF+kxIEjJtnC/42VDTWHcwcPY3JNa2c3W09wU7mtAKyMSig0Cnx
+LnBbSHRDlL5ByQwcVoB7mF4jW54Xdn//1JsMD3ALJTRnIrZ4D2yPd8MsXd2MyPU
6RRTqZ3gVIz4GMhfLb9vxdkqog/LfOUx8eGKyFjFUSXDNWUEnP0AFMhZWPNTszBk
ZT1Rtgpz1B1Wt0hl1e0xUWtX2f51XN1g1qmy0LNAJVU=
`pragma protect end_protected
