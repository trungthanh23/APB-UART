`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nNTtbuuONAvF53X10unN/GCXeH85FzCs9xceq1oPp9Dn5oQbg4TVzUgmQQbP4qXW
4SQOpJ+k8glgjj3yp2juGMmbChHP8MXQPZ6L4LRXjZoo5bzMc9ZWaiS3zo19BBE/
W4gmWHrpIqR3A+m4yRnGU0hRL/tWbPs8tFTZsRv7qYNefCCZCkzFKx1spmEO6MpL
Yu99Ja7nhyoWz5o1j90eCI5Af4Jot/Lv4Bre/Xa/Z8i1wzvvMdALNbVcIQKkXTvI
jKzWNzooBidRWRXev3gMCKjt8r7xQuVePwHnAFLQvFNGDvv5K8yS0oetxZgCtOPE
9Ys3JX7HItvh/ROOA5OYeQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3744 )
`pragma protect data_block
ITqZF8N441apjtu+6a4xq00Fj+k93wr7+DlBic1xCnjeu1xxz8FOCloqe5PGB98R
0HM8CVzlvLz6mn5eNeVey0WVvMSNbTrsmQ78FLAshWa1yP1TLxzrJz8KxBLA5uO4
DosisWFC90Hp6vtilgp8vRZQdfvwQy4ZThM7hzNmi7ElT2UWEbon9DYDQqstTNPL
UFNq+bUilPm7aFgxN64DguyYuDp2Asxag7EJj/ukrNwn/4nhF/vQhdK4Y6DUd2kj
KdsFPyyr56jUrCzaurGODeS9KBzXdrUMZByWAMommLrixf2v2PVxDLZV2JpD1GXa
4uYPpoDpj7l+s5xalaejNbv/FzkuoOgt4AdQfO9rk6AWTXTjHEoo0JotXoAvtjqm
oMgmRpF1UkxGYs+ykQg8y7BSKcOb1j1qgBCxj308v6JrKJ7dD3YRffEdykxKJoSx
ubcCoq9WuRi3h735u95m2VgyNR6P+vFQruK9N3KAXR1kwZrUKWzlOGwE3iu17cEj
YNA3yoDJi/ojfMY4avmvnGE8bPXLWtXfNZnul1Xw58pi99A0M2BmTFsIKcNyApmr
EAImABaLjch71XGnDWhEu+CoZ+nfGHxnvIReI9w9L2pY3iIqjwGnmTN94W2J67xQ
kZzfc4RoSqHFvYiHa8RL3fg57x6EuVke5kn8cBsS5dRbmDv3l3FW4I+SPEAUijHi
OrdT2aswJP0wtprtg0Dlh/PpOpJD13kvtwVKZehMwmdgNzkxUrMNerWXaiKvFEwI
2zGqmQ4xXMNl/obGeLTWwY+iWslS+HIiOUGHv1z7QXKwUu5V4jIxLCp45nC6udF2
/ueiMwO3Rl1gTyNKsG0aHH8D5oOtZbjAs6Sa/wRCSxdb3TGE5rM/PzLWNKBIs0ec
9sNehtw8bQsxNBMf1yEppX4hFpsXhNoGSSAbM8ksBS3/q/K+8IatV5CJvPbJ2baR
80nJJKQn9/8+vU6RY6Slv54N9QHdBf9zvavYPvdcoZFSUwjAWMx++DKfYMpqBuKF
q0i0yjBStTdfNm7Azs6BMurePzmAFQlWUoDcA7x6mY1uw4FkUVJGMcnKx4Czwz+a
LQkTDlyvHfVqwXteFtJjXUK22dYrRcHtr149G04LexiwW7twYsA6SHMwpc6YMTRa
seTCY5FYVT5BrDBmp5nT56RU7Xj2qbbDoZHkz2o9Hc2QP7m/JvrdWhULTfyGBvGo
Jr+eYQIzx8CnOXZky6IgcJ/e7ugP9Cy/VBa15jvevDw/TWUXBj8sM3PY/yL9a0Kc
uqoD5em/Yzx4oNobjflfmEDyCmR6DjTFi4xcxsWT6OcrlgmkFNWIKVCxF/eBZfZ/
8h1zI2nUTpQn0rZayFbDT/rqGrelxR2qbSh+xbZsPauPItGHaW2eAtRy1rLm0Wa8
y+avWNgVqFclDX8LncaEQIIjx1fu3QC+GmC6nrDUZxj/BivxuHUj06lPLNtqeCR+
3hXNnwQreXvk5glsYwtkWdtwUv46gN6puy2kL2IEFTnXA1uGgyy/TYRgKiv7nHE3
e855EoUBYZWRq9AzalKTxb43RTBnXCyjE7Dh2ANaeXz+0vU2ks9l8UW7TSmxYR6u
p6D1x1zSVFtSSoHcs+Gv3//j6wvy0ZQAa82e4K3Zmi2HmHMkfmWtYdlN3W6y5TzN
qBDw2vX3fN11pgz2b5/fqdgD6La2Xteyrtrv2uAlp1UeZ40jMy+GIafG85O0Uwt5
sKiDCBg3oLyDIg9HszVZRAfduAvSeDRpsQziqT+YTerbG4OZpnziM25hHFh9kkvB
CZ4ORAJicWtOispjkzw/4Eu0tAqiq3jZOuVIMIRzY99i7bFNGQPymSmZVoByJKuk
XPUehsSP+2UE4uEfZekPwchhHUqrwUO75aWpItOx68+yZwfiuSkupQ1E6LwT7Cl2
Bxr8szxEfeVnBdmDsDCzwXBoWo1hj1m/4B3iuwXh6k/VRwVtL22UU5p2s7gF4qrP
0J5Cq2Q7Ji1rFtZNFOqTeBe8YZNyLnj55BKY5/yoJFDqjylIL8N32O5/USvEHkWL
iFs4mb5+0x5KMGz5c9kc99HdM+tE3b+VgISPZW+RkB2Egopfzs0bLpcVFPRu/wUq
rlc+Etc66T/GXsSMDN+5uWv6AnfKHejT3fwJXao7t8xq1EL3char0WWiYAip9z1F
tKh5aT6+LFCh5d3/VBeqQpdbmUqMgQ/+lN/HDS5miYzIaT+ngxylrizoaMWv1yPI
LHF5Gkwd/faVTFDdVUGssKhCYzL508Rrax95pZhmS0NCVHhHt5Syk+h8gT9GpQd6
qpwgZseVnfsPJOJJQ1OpxhAus0plpGBNaaQR8j2cGLWqdI4IJQRxxrqIJt2YBMDc
4Ee2OOfh+SBAKrWNTSlrLfjpsFQQV9MteO0XhE3KmWneDK7LmPkYAfQUDnywvNRv
P/bFPSSTCydqUx+dQ7Yl2xi4PVNIN3wSGghqpmVGosOoGaS2KueHWIsq1Dt2gXOO
AQeoHzLC4pRLSMcRzLVonkueVLBQr93jAs4yRNzCicoBk9W2nAQPFID5MG5QRyA2
JEWMRwcZcz+3JpvIgSINd2o13QU3qKd3Aze9lIFtxPUe17hjrcZctuSmHb1U1ZgS
EvBYy/SFEY/Sliu1R7UbA5V1XhnyDNu+LhMl/Dt48FWI8TeYO6ij97L/N2RMyXdf
eGx7rWXQx+LVE8X3ew7JPcllyKAkdrcV12rqW2Cy2ycpwQvoDOI/sTBkfxCfXJQj
9PzWokDhE0y3Hil5SNB0MKNah7ZBX4Q/fOCBoSwl7BeBYhxCp/nPCB28tL70fIXx
aJ+j1YviKeBWC2exSCELojBnxRYSIU77oob4DWDL4p7deVGgZfdwD7LknM9jAb8O
W+JslGeinEJPN+fgIXVxCpJ4LfoADjPLDqnW6KYAMEgXD3PJwgnFWbgTMvSsiRtn
CiZBfX998Dq8nQEcxQvi2YcddKFCmnaLCrHoJmCb8YYInPx0qWoxEeLyEkoEWQbz
wqIKM+Sd1vIUWuOmGnsgGjQwnsGWwMSTu7OG0n6j/t+AwRqRB9uQmsLyL9jJN0nM
dvgxWdcPfjTNWw6OSjYaJd0NKv7wmOg4LrOQ40hpIk6//iWIBH/muc1sF1oN8Dxh
FkeX5dlWrsabGvz+RttbQspQM53Gs1rb/JVyWaciiykyRblWgD7lBhCY+RpkTLFO
t6ZX5cbtqv2YiQOp3HmjMCTQTASZz1MT9YctDxUNgqVSLCJpoOe0n/6c9rm+hwIg
5w0rdhU0CMreimZPQ5Mo9a7pd/YosTecWYLMQ4p9F6smL4P6VOd4eWfeOKmRjMpE
DY0BgWamSw2gC1tHcgxSvnElwWjO+5gpUzGTik6F44nPe14zhzXN/htvsb3k+K/y
EXtBqWmp52BDmeFby/3/1GY4x7wMcFG3i2GgD0VUqrHh1AwbJYdWBp3kAVENiI/A
bzuiO27iDjsLFky2XsnZ2rudg44iH3XQexVeMXoggr6IdSM467vpFHgX9RQtELh6
qPvxmR+/8Gdjb7N36L6tMF/xSxab2oxbiv6m53gcetpxaot0M32vyhC0dlXlaZdp
8Ja2s38aAOdnlQGw6+Dj6/9D3Blq65RlJc2v8DNnJYhev+OSZuZS8raofasn6J4x
ihijYeDGcufWBNLHMR5NqY+Iud2y7yL65iis1oKcaU4DFxwQFsXujbEILzPVJRTf
3B5PPKLP6g96vc9yC97IloONXfMVbqJyNeto6T8QQ3m0Sa3ko8urNLzu+M4SrmiP
hKJuLFekV1Qy/cPu2yZuBsXAVK0+VIXN6j3e3p0/lMTQjpIR6o4NFo8rs0N+Bc9v
ofuZcLyiZKXNzuSncBTWDshW6N4Bzx+ix/OB6v6aZSpHz44ilICJy9R31xgsfy3q
CnArMz4ZAtvyckv/wdqxh9PAULDhTO8LNzFMsg/zjpdrf7jHdM6WgZv4QfO895Wd
XUdI+pTjVwAf2IseIwEk3UkOgl4V5l/8OJeOxCWhwHPqNslF+lZFf4GWu/20nhrM
kX8+k5qn4yr+DmiG/CLN+2aCJBgyO+44gT8XU4R8fiec0/1D3IsX4XAC2Csb1ZrO
ZFzBPIz+hIGEu9plXLJaxH2wZ+HdU9Jxn+2eNAdTbWPy8EuX6R6PrnpaYKGo/RBl
wxUd4imm5FcpH6H8hlwfZ7zN3dxtJKEH+WPvX1zYkwrHcCABGd9fqTGEgap2xUxa
PGOrbmcAchWQAO0l+V0bsTYFcrMabiwPIEH+PBA/7d1Np1MVSAHOz13kR+Eg88If
YjvSnSe2ZxdkhgE6Hjwu46AmVU4MO61kbkP+KjNgT9uuS1F7Shx9+ULT6ETpkvtg
Q9e56nziLYtFl/PGQYW26H8PiXmJ3CZU5HWrijgf/aoJvRYnDeKLNCxcnrIlUC2m
ygcZQTLbKLsxqZQcnh+lVBvvI1vcbz8mFBVwU5G1/7Fq5QvKFlgncG9zeGtoQNbg
hUPzn1BTHcUWJ84OGj6Pp1wTv29gZlfg8Q9EmAW7cp6SzykVBA/zNWNDHdYI/foo
GwRJhyweySqv0e4DEsN5Cq9fZ0tMijlQUTE08UaMs4TsHQJcWUM7yJPJIJocDyKD
8CTtK50t2s6UgLxiXUsyjJZDtbScVVeajTTPLFa9B6dIzUk+VfbE9QPtOLYxssFp
b3zOGRY8wrDwPNfTrUgrnTZEinJAy9mgTylj/Hdphgru6bfP2MIFmyXAaxitgfOD
LnCg5gQfvN8Q0P0IK9NtVsDPrjbOkhtnpGyjeN71ArXELc+NBLF0qzahFzXL/l1u
bIkCmhhosgcIPtYJR5lfidHVYYNahGkleglheHCgQiRqrjFH7ni1qCsRsOcE2nB9
TK48L9qczsPSAqgg5YuJJv/fBzZl/Mbp2ier1x4w9PH0G61ugM/3eItfUgS4ZMhq
FQHE3/qs86NqiceMX4EYbc7YczXIpyZItl6Bs9T6sfAv45RqWGCM5/PKQKTB+vY5
`pragma protect end_protected
