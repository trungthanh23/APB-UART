`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
i2qqyfMVyIylEbQZa5ocQ3tOEI2qaMGutQaBAJv0p4mC0RP8SBWmTWXmymXT4TWR
E20OyJxvFK5EOySYLtmPmJJDb4D29e367rLPL6pEL/AdVK9x0/Ow4BWdqx6FpsL2
cfDmDRQVJ6YoeXKfo5AZXGdE5pz2ChZimXrxJ0xtjzNs/R4M8a5PP1j2mlWcGSmr
rHE0wIwzq5eNfsBXYPHybHmrIar0VM6tgEnvtvgz4p2AW78e3oyXJUlcQRV6sxnN
/L2bPxhZC/5hGgBGl4EpYiic0dEJuR4vdbYwZRGrcJExjrXKGhD+c6gsGBLYfiP8
CcelXT7OyCB/PGKhfC5jWA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1696 )
`pragma protect data_block
0Y4QwkJf95Xq8AY1wgcKk9UllKV7i2PkzH8Y2NtC/oVNSEo9IKuOW+yL6zTw7Gwo
ijyAFpVpJRWGnNaD7AS04g8ROsPyP8c3jCfWXBBdIMQiAGtEpXGY5tF3J+4A2Kfy
/STHk2fw0/mDhIA0VlcDNfnXbXXZGcvIyGGCVH7tlEskZ9XhUn+tsXuMfNtrzgRg
45kjQWA2L6bbHnJD0iWzPH3HHszgqaih3U0AMLf8XUL9F8zob68oRPFUGNeYTZSD
KBYTrDxbZbhosLgJwSCqYc3Dd0RTTaK+49XYlp0KStdqBzeVh6vkAbobcSeCXZdF
dltSvQlg/gKl9oXAu1z0kBsmYX8aBlqAcxOvxKQmc6vJB5KZEoR13+NVMnmMKcVi
p/fM0JrlRALyWGoSGyIgDTKKP93vT3Lc4IfhFYlDzqg3rKehaZC7mbIZ6rqPVzIy
qoPhLzFT8YytNv45XWdWwlvgX4CvxyVvFCX30fubWbjotV56uT3gGkuCdG8SgY80
0mlrJxNz+p45u+1o5dcnjGnGTg5YVRIuskayFsgs8IqgH2BIsCQVqzveqx4b973q
WV9O7APrQCzNgEtJLkjQu1+9rEbTts77Fxi0/CaQeMv/DuS0TitLCguSlpXNWHCF
HvbugG9xHpIDYWyqJdrFl83Uv4i8DvNMCjHF1ofMed4rfx64+YqWxjJH2v+PNo1r
B8ULuepAli0pvDxaLLXRD2n9U6Ogqy9r96Tme3nIHVgCLVLMI7VWNrN8iWVfT6f4
Vugj6UMQTYRL9zQaRDVSMIHcA8/gKhiphpJiE9HZtTX8wa6409eeK9pW8cSg9jUE
zud0JwBv/W3KqtQiYNLXQ8bjpD1jhRZfU3UvU9wt6KcnG3d49e5VtFYnarVtAXfg
KS27/CS82I65gZwcO/WZ1GhkjMPc5tRiHjWLZfJLhWtT5WEIcu6b3eX5xgCizJQr
XtMaaguWLrIi6K0ZeczCyw4hd1fgR/7p5oeG7PdREiw/H/Cf3JMVmCUy6THvhSmu
aZycsUYJPFj78Uhu3C/KEXnijlwacUWrfGAVIi79vJRIR7y/urLLREf7KZfWddGL
BJvUQ6BwtHQA2IDD//JWVpC6KBy/RcPLOZHr9rFg6xFH8f/kouhugExlt9IVUNTL
jSiS1bwnx+ZNldr/wwgm18eyPJo3BQXbLDMr1DKPD4fUtSXRPfQ6+9jv4KwdfS1p
z9yUEK/nA2keamZQQzqBvATHBoVNiCyzwwvE5sPbKaW2PLBJb+om8WL8KlG9kl73
+dduJTfnE4TI3iT7svkkaftQGXAY9Puc41YQVTKLaOeWcGBYgb/UUInjy2SLWFMH
WMnhqFe5raqxql3dGNc0XXQbUCEn3pAwz3vuDg7sKqAgHFa3cBwgCL3wt9l5Xrgp
ghRDoEIoI063W+xRVGA349eaA0Ns8UuQsBy9ahONvxH81aDwkX3HnSXjbmDubXNS
QOteuTcUrM+WlTkQ+5cqzoxR2BvQfq1+jfoE8OTWZXDd56vPn46/TQPdAgtsLg4z
aZZhlj6oDxMzxmNuDtjsAfIqISOWdYE1pcOoq337B8rvn+fcqcqQXw/S8OvfNfD/
U7Pq8HUKX9s2Xg+tt4FsVdn7/MIDGkoGmEbbf8VTfPZcxVmah2L8ek+P9veRgYZl
BKukhVj8BjFV3sG1rhXzmuVHAuQNmtTBdRro87+qNo5xY9JS7r/n5Q5zH+N9r0Mo
V1tCBxBBatTU74+t9nVXaGulGYHt17CeM9lb4lL8hxyrs8a4DzmAx6O8t6dWIr6O
NbQGrQfBrQeWHyTkGGJ5ZI8ry6a0q2IaJi/LwHvLoioIi/U3U+BxriyQZSycDzXZ
1FfE6gXPespRyf3eCGTIFkUOmqzHQg95/1ln65vtoomPpg/LxeSIsDsvQujxoeZm
9VvmzxdocQZI9ybsRQtWssiUc1jU8nyP5QSYR95i0FfYKRWWsJXV8gMluSDZlDY+
oA8oapIqixEy9XWKPRJjOxojyGY94o70xWPd7oi17F6xzMbvxbrY35stVp1gpHgH
w8DwimAPAfdsc+yX612436d0AecUVljht6Yj1pYacTz+xLZM1+NKn3qDMBgLDVpS
wYEEGg9IX7E1ouPt6ht69QNfsOb74qdjR9LNXPFaU49aExzkHO8EpPT6ILE6w3VG
M2FVduPGEUndbnxaOgeXxkTaG2kt5tP7TcXriNdEWnnUSTTWGjoYekSrV34yh6ru
iRqcekP2Cf9G0eA685JOIg==
`pragma protect end_protected
