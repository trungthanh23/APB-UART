`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FvDzw1OjBIsNkmXUZNWalecJ9puhDQ7JeE6uYilXqLXPPjQxuLc6hHnDF8vKCmF0
UZ7rMApv3nX3i35TQSo4LGnuZV31d8f1cQ+f7BHRHmUchH0KLcRyObrWwqknY9/R
B5dBawYq0jUbNb8uUHOPhfbjmBG/1GKl5dn/45YkY3UGx+f4uU0/eoqXUWit2qg9
8KOOB9W44aJbCElKCDDs9mhCExtF9jnfAgITsP9NUKNcxZH7ftiS1Ih3fqCDkaWN
O9HjwN+xCvswovYemT7v0sKjqnLNQxIqzjmd2M0HZcORCZshjMYDpJtm1EDv/JD/
z6n92svd4eLET5+GCeD/vA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4144 )
`pragma protect data_block
cRgp+qf74Um8QinTW3mIO4+4hQnJzhUiABMVus/BQNDwGI0hFG7sN/xtj8I1YbxO
z8HQ0F6Y1pEXCKHPnPZxSnyletMwl0OcBaD1ICX5CDWIRh4gA8TCaXuPud4RZxbj
NlBYwa4r9sZifZZX0csKqSolDFF8AWSWfBP7U3MrKPwvRBkAf+9oxLSR1Rm642pA
cacngbJ2vogcIb3bBtE+9jE5SK82KBzVObqZzp31GpKyckoFRznMs44O9jVBz73H
+QkeJoGtk0sTsZ4lqbFfoVpsUEthpmhfIMTE5q+Xpz9hiczYikkA5RiMvR0Y1o/N
RDO7imnGSG378xfsTJFZuSD4lF3SXj/deKGwa4f3lpNa1CS8iv/L8oOeF8kCeZj5
lzbceVRIUmoO7+/N3A4OaimRqBZakNsnRmdrXh7g1XH9h6wfgJMZeZzfP/hB76WC
S1vRDzF6cvrtQ0kBejQcwj5b7PLthzRO4J50Gn5svpdeXBIiZETHdhIVZzcZ1v3E
iZkdwKwKZebnzencl8Ga0b1BF8vonkXyKoBnGc/3+1wE7hHjBqlEu4S33eV9Lqmo
cPUKjUepDhpDo2Dun0qpNEzT9pVkf0PuODyfIu4yS/bcVT53wdJKzSJC+jRaQeGI
bYOl8x1Yi0TUwwW8LOPCHPBFmTvV4RsDv8ElrJ4sAoomfSsgZgZYo3xVJuyouak6
p2eZIx0hV+6c9NKPAfWsAq/vbybmYDzmAMOTMi2uCh3xg5cz7LBDhPnLrG1ONDMd
DMnn0KZPDUnNxCjXEANgL3ZtW1rtyBFrDEgU8SOiJdzHSJezvpVT1fTNJrareABL
yFDKbaBSHa149GYtbC4JuLqyB+cKeSwxqzSrubPRPF5U89vq84ViLE1ZcoGsCi+8
UhVGveLJF9j9DJDMAz55XdHhJBW8245OV5aMfse7x7reFPl++OdDRc/e1Zj62fqs
cJxPa7AeqEYrBlagAmsDuZfbN8qp91r7I1kFRa1BfhZlBz39uCg9BFdBUySRdt9H
DNAXxeUs3w6OAck7nm1R+NU7Dtn9o/KBUYJEiah0bMIo+WeAuxUXrTooy6DdnqoP
0LIPp1AKyHsZNnMs6mf5ffSsn3PWcKVFNzmtCeGTt5BuILlTzTSHqtYG9Ts8GvbX
Fgg6bL/IpDOojonOoU2jzrYp2aTZjXlwle2GuiKYQbMxTsyen8rRKu0itWTq9XAc
zHva+ouGzQpr+h7ZlRRzvXhV/4rOnHyi8l/k0qk9tK171BAEMuvMGaQ2dTGxjdfD
X7xxNkZEOSbQFPXRuUQUCbcycIIlPEaxz1H0sumxVXDcBRz0MybUkyeIlNM0DxGd
+/PSpvzCG+91syn/lufAseHWaGDNddtrqf9CfHWUIQhq4lSMKnxucl1qAiCOsYKm
IP0FG9P75dx2LpMimo8OUSOssq5VzpPNJSoyJB4nHbBsktjW8H/VYKfFQR7AfRdO
auwUpt4bq4eILte7XUozbk0lPjziGZugy6evyQyqYiq878XdAL8s0eQbPQsTviJc
Ud4DolMtkpS0/MjZjNsR+nwAXbmcfTt4oHQ5ezpHTrV6u6wn/TeIBv99Ll5+u+s2
AZOJMNBF0WXH+J3bdfTUeh0CATKSdLBiK07F/7+5qww/tBH7JICejgjFXQWlpJXn
QBg5V6SH3qioQXLDFlXEoK0wdWLW73X5U9w9gUldG606fqLduwOrf9c3HvvYhyfb
vZAtQOusJF7s03RiQ7RKcqvuOz5fAaPtcKwBm5Ho/ofV7rh0cFFpliF8Y2Hqngvd
Loqb7BKI/AVTntG496Fz3Gk1kDBMw/QbWUfkmGjHcCPo9ikF86ed1ttNy/jGPbig
apnb0LicPS9584LzONXLNX/eVoLqTJe11Bl3X5GjTXALTDq5xPvSbg0BceQqMb37
DTlwc2F6vLzD9AzAxXzEAlJ87++KA6PXfNiPhA16uh4r40YsbxvuW1tmKzHh1/oU
41ro7Bho5xa1q0R6nXl+YmbhF4X5obSU10NIMuRF4BOiECTfK9XFAYHrgkjlwxUp
sfXP2yyvovtISbaCJsR2Z3N5Fwz2y/CtXXUMkf0WpzWs+v4k3Vzy5htlFLrg8E/Z
Qt3dfQES0hUanhboCGgdmFnfaclWUkTS80PN7Zb1BRHR/j9iFiHgXvACE8muqpc+
UUGGsMwXS1yx5MWprih2BTowD1UJ5qsYBAthOD6bXQctGEblcy4OTDfD0on1usC2
Iyy3pSAo8/wvOPqVsIWczOAnWCLskfCUVL/Jl5l/F2otQjLhpjRynj4n9Mrx6b/l
fqBNabK/ZM1JGCe7YC9z2ZAVo4pl+T94p+RZWDg3XmjECTkB24Gq4XXYr7EHJUUv
5e7+5K8q8pF5/JF1EFsRT0KifBfadvt4imEVnqB4BHyTiP8e+PytirtdgXY/sV9L
1QPC27SyV6wKCLwdoylewsuaY4TJkd2IXyAo6R/PHvLp28Gno31KgaJMDzAMfICz
DEalNT3VlX7yIWfLUhAWXG1Ros2rytVyyfIKMWCcEx1o4HloOBgXjes+BwGR9Kg9
9/SUum+5o7/X+Fq7Cp6iCB2FbloSATF41I/cKShKLOgj/4WBApQ7i6r08wnHLCLD
wo/z9JG6G0gamik8dwzOLd1nKTHS/ELRUuKeOv9daLSkR8xI4EyuM1aVoioiHYW2
IkIqt6ykU14WxHJXNQpTU7JPtngWweEvdQ06GGJs7uetycfzGT5BD0VuiNlVT5St
zLrOzekwpRmzvqFr2RHDH1xs/6lR9Cfwsge1MzcdPA3BpcNhRgYnW/12+Wh6vPzL
74pczDcei3rYCdMnq7n9AsOoIIaDfwU2Fijp5DkyrDW7269LyKQ4lVQbpFmT4zkE
MZ2HLugvgN2XrvWXpOCGpmztnna4ZUrKzIno2EY9Q21ltnOn2DylqRFy38qG8NAN
+A2UsoGxJD3/+LLSctJE32/R6lvVpv4/bpwlnkNMULdLWh3LRZHe4+Pn3M74XoIR
aAsYsI0zQlGLocIGG2isC2g8X9fOmIh5ZqYPWu9v4Z+iPr7+ItcR59U1FoJdz0tc
jIijwawS21ht85LjW0cEUw3lR5qt1CTJJxpthuF7b+ntAVoIjE6FmDs5iBa6NONF
uDd/stLoFO/rLZ8cnzi/bp/5IL5/Yyw+Z+z+k0XH4q7yYUORnSt/CLn/IGf5EE1l
K/qsSK+GVJDks3f2mnpFc/fE66wVKd/u1Td9hZe7qb8CdCn8mPS0zPOaeSO2/wgK
NYfNXoVDDdFMf9OTQC6O/71H0fR4egZZQ+avxDUYTi4m2eeiExjjdAvGTjkojeV9
UHm9lPQxpK4YE7pJhFN8xPBFXiIwdfvu0pZKTRo/HktEQO0zqiDHurJCLrhby1/+
bu/l3LEHaNFFzlytp8b2hes5DsPfQVR1atkN4G4VzlZ0nTQxSRmW0cZ7o5dxXLv/
5JtD+qjffHsPcQu8IQznRhrJx8lrls2EdotikKMKZXiJiPYEEXAubKPcO76yoG67
j/VfjBnDkC4jMabVXpQIGylUyt0m4x7weSI146cn3TUM5wG5DWZwhfqyOKWmF4vm
nKa+UzO+Qw4h6alDbP1ePMehDcv9tIuUO+Ewa01oIVMEIdHHC90P90MxuFbTKEQ1
xaicKZWyuEK0wkyWdH3/tkEgIcWYQTade9RifbTcJeHGRUYcGSJvkwBk52PtUD78
fLF8rsRGl/sZ1Np5dcX23wqVV8NJ56sVskQDjcGQshv3ybOEfKMARe94EL3hp7Dj
xS8hgM4KoUPAd8r19ZRkC5FNKNlGJr+GvkttI2NieQ2ON76tuLqhZQe9amdK0Rzf
rfXomGFwfyfzd3DCTkP65hQW0o6eHBxQROWNEkNvtdFDK/ROlelUj1YwMbLBpE3R
9N0uoKl/KxAspyONZ8T2zp0tLeGuWbrdz2ZqykzvVJ9GHOIy6mDB3P/SGV/3s1Fk
3wH5WD60YqEmIv9A1G1ptxPoxRCEMGomRd93Qgw6nE1JkhVivz3A6nUuph5vsRgg
niv2yWZMI+Kxs0AiHCS3FqRqtFqjDRrSMiS46pU8+u6ck0NIUOf2S4BbTca0AAxc
eUxLZ0T3jxEbXXtpJ863bSaZEOkL/Inj4Sb79q70JO9ICeMv/rrhmRor7MJOSEmY
cdi7TIHi9Fl2nxQ3I0UE+wlVfoDV4CrhovLivw9uurVpDnwtIcGvvLxOvxV68aNb
V1z2lVDngb4iYEmt4gNpQw4i9kkrKh6d/zKzXoPbVLKIpWFFFWlwSDZrDEWSWIU1
ENnFeGhMFlk0Yf8S9dp4WiSXlI9TA27w4YTPXaZ6XSn1iPB+xCg28rW6I/lv9ifx
IQz6CLSCUhuwexQWVFsZ0SNohl5f0LhaF0kQjPd1n6hoxxsUql1Ck0mhnUZc1EAZ
MrhRHTlrvwfRPS/B4VOTor7Tm7DEjTLq9+TMGRjL7AvK697SUkg7mwLxwmqT6vdp
Tm1RaVjJrqe+eIEOJ2hkg21GmUWnAQFbgDJGyx2WPhjjhLpL/fvp8LcoUJQdWops
kqoTcoAUghmGrA72BTmfgWd94e01692IeuJMpgcCw9LqUtw7KYrb759dX8WcepKA
our7Fvr6Uns5lPj3x9PW2eLiopNqrIUiUqSItUbfq8ZZsCz+mPP6SdLuTZ3qFZcX
sb5nMpyWgQazC3/H7l3WTkdWh6ZBPtP2BOI91aGc1O66srLKUBHiTjfztdDx/YcE
DXBa/LjXiL/YM6leIXeTrZs2PQBQvg6pqlIWcPlgok1HxBPBHFuv7wy3sBKUJyNc
We3bA3bkRX3h3ng4A+YbaW7HhI+6ITvhVcjm/YFNKjexEm8WEomnAwLlVmdWlYP2
KaWmKDXEIVDFwcLMpcT3aEtU6poAYZQbNGnj24VDmIfeTg7ZRrZC2l5EfLTigPIe
3tPRwyenWxyuUTxjdoEMWNzW7Cg3MJwEj1CeB4JSw8VBQe+5gHEHpNWetwrbxsk+
fN3z2oMF7YCEOAUMqVzClk6KJU/CT7ghVz2IEC7zWtPhXzwg+0VOHQvzdz+ruxWa
zNoaXv+ZsYPEsj908WYSn9+2tXejNEazkx/8voegDORhijk0wJoBuNkvsxlKomv0
TUyGYE8KbFtzfXtK1QBVQQY/Wxv4Dm6Bh1TDmfA5BPMJS5xM04A8mSrDw6DG1MaQ
CJ5Jt+2Re7O7UrmgLNabvuGXx825pxbxQ9a6XptjR5G6WmLlsFNgSdBHi+2Cp7qy
arI9/7fpfcmkxunFZ6EKjeFVhJZXaDOi65UCMLyxLAZv1cqhgAJn+b1dNMsnYiR5
fVGBnNt0E0Gwr9iB7vCINuA4XmUN+TkjVacl33rA29wMYItrN+SavtuCvv6yOrRA
Vs3EKpX3bzevp65TAxV58iWVY4KBTk3u5DGhUVMgQsNlbxIK1T+sVf0DwkWydKP/
iG+UompRgEVOJId24Zbs7y9sUVQtbu07waOgXyXFoqJQxWWZxCvFCdocGChkuQ+C
8xij/A5OuU+D4ftPkMiEAw==
`pragma protect end_protected
