`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
DyjqzVWi8pahR4DgFTYpGUfYx6B6r/74/Diud30bDx5ewKF8wb8gOoLAwuP5Pjhe
BCW87T5s58tTVQZSb7Qg9a+eAO5bn2tfkvac0BpdJ1IXtIY1emA7nB/uZ/69iKqp
6zgJqyi7Ssp8dkk9wnxB8jYreYtJjgloMk87M9mAz48yXebpQpNw/l9k7alohIrp
kkgDaQ4UNXKyKA2R0Q/WZDehe3VbXz6Rc2Z9qEp9f3szU9oC7clPMnLSjhvhY4Aq
CnQfC9EXX8454bmltLAMXNcbruwtLkkYDdIzgyQmQWR+48zuziQ3pe3w3VDxUUzp
pjONgfwWkYaKzzfeuy9ixw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6640 )
`pragma protect data_block
Bk9Iizvv2HoYLp+pkhcX0iit2XBwHgHtbLrPp1NZQiiuqytCdoddyk/p/VtrFtIi
0cBP+WdR8WelT42PvDBIlkOF6Up5gCs478K+HV9ysb4QEpXqDYNbpk+yL5LiJnB9
2z0ofNuN5JQH5j+xxE6iqwXRn/M2dM3wDU0p+//agFh3PHXTJDhbHzzB/L3tItkj
rtWIRTlu83N7g9ZRgA+wFCWksqjZ/AXrLOBeTXdDDooJX5mMX9S0O1hsR+H92gTA
BGcFD0BvFUmgiqVaFRkqaLuXWpTj3TxNskkg7KnrhRgzb1KIX9tNgU+UrUWDToY8
V9OWFzEfQezndHDYmqNu1KKunn45Vuslt6FT9ntQJlTALIcoC0CbLgBi7NPYBfRz
TkrN8On3a38R+iLnR7YD048MNEqF/nsfxzyCk7WFhtlumnSYZjVhTOH8xTp6pVtU
rwgMom/mpsL0mKEvjhPZGba2yP/s6Zif6C/sb0/bSlJdIkgEJXoxEZuqkNS8beaE
MtL1dLaYS1Wz2LM4RSSDx8g2joriqUOCBQrTqY7q+TYeTaqJsOLbR9lP815GeO3O
YuWTFBkzAt8KLn3TfR3bMqBjZYjDLLmpNtUZnAPpy/sGGlEsmiIH4iqz0XrSLboM
DhC19WgKwvbNRXaFuVqVbjlWwJjLGNXpnfTDp82ML2yXVnwXQiIb7JE3lb16N5lC
I5X67oJ8o9zGZLu3K3M9h7bWfrag/SRWpUodDHHLxice2xmjhMJVzqHcDph3aP/s
QqotLcIth43TWPpWwi8MUJBu71Bz6AEAFVVaP8o+Kik4ku0PWmEVRDkcZFAI6VCf
D+yCWbP2ILcmYdbBuTaAQWcRF4Dk7W94s5ROyPYPtshEa505EmGiPcpdKM3+UqCg
i34T3QZiFOKvLNSEq9ndpR/0huoq+zMFdPiMq8Db59BBSzV/5f8O1TLJB9T3clre
xhOop6gObeU3SUtPv/9VKbbFziivxS3nRfDOizjJ0vjn+UTjmstkHIEfbM821nXh
GsvPQ1pe1fqNncRZRxI24b95SGrNfA4V+yU3PCmXh7t/+sicQDAuTafQLfZKuDRg
B+gtHQqhzzcYvOQq/HGZlg3OJ47ijaPXlSZY3hosti7+K97IGb1ntuMAaxKWdOJZ
/J1LwhgbxS9kqyxQAx8vDT1W4tT7E5ibl8m1cLbkuTIgeb1bBxNA167gBPSS7pWV
UWrEeZMS902oPpP3UPlwN+wbvORysnHn/wdFKCFI636oDVqmPnE1igl9NeRtPpNS
Fwzmfmd3wjFdMz54tWnhktd6S8xJLmcPnInFcuZtknj/SMbE5gCRlnO9UmSIJmSA
sogmJnWBtidwaaoW9fKuZyRq8b5CpmeECpk72ryQTkxAELDOcmpb5QYfbb6sK3+2
3t/xJ6/8ICfYk1CiNNQij9GXCSPLBuBe4gLYHOtO5O1PatrQSMTSrh5NTyCdgOth
Itd2saGFG2tK9hEprd1sYalSK/2NWh2FYr47pCe6fraVWR+yiXpjJaWXVFCdSYaz
wrgNlI8P3G5BQTDgcdpTb1mUEDhKbxYYS5ProC8SjBLSW1nAxJmEhHE6C2ZNZsMG
F/snopPo9+aq3o2lwIfQPgLTpXaMHw2m8tMl7mUlAGGJkkzelrkXLmJxaEkHLOGA
OMQfCKmJnF1Ks0UVH1Flq0LTgQ4ZPyWSuOZuGeVb5DL+0SNutMDn5kE+hcxfJ1I1
NohuDq5uRXwpAzbAu1GEVIwm4cIThZZ/9JGwBUBmlS3RKaz6d6KEnYqbGtUH+C3d
5lC93QlS5Rvfi4lUYtiNYnTJrlQ575eyDeEK5HalcZXQMwv+lPXOW1pjxdsmqKQh
UUPcOLOmhV6UNhGq6OJq6cKhvEk02QdH1OxEGICtnF9qNrZnLO8eYxO8tjXXNMps
XQU8Cx+Qwlx0p0j3/I0L9cBjrE8LG6zKaRyQci1LCm87A5xcwiptVc66SnaBV4un
Zx2kO5uvp+flfXJlBYDpifPsbwF6/r6sHLP6OxVDB2e03QunPx35EFRPa2T4+DsS
bE4saOCUAh/QZRtz58wcKYcFlK6QXxC9tw1S/b8udbE4TRhKL6aTYZNbzhQdJr+C
09SRfsr+8beys7/uA2XPabplRO/YssfFFHE0lNJFQf8KQZA1WydQ42bnU4WH3W16
BG5bkkQZ53jFmUMW+IsozgY+iLaLgwRnFhVhsB1cRyHkYQXmy3kdaJLLWcvZZVon
jra/PouMwjARCt+Ms03IY6qXuuuk7GD4G1ruNYn5Ik/PrBQKfELFAN8yR+lVzrQy
lwnhM/qdkN+ppP0dZpA0koH6RYzYo1cMJ1GBtfk4BPjudwC6GRhw6cWtWcUAk4wV
81V9GlHJ0E38iVzlvVowq0QI0+qvY31Hz53lcUXAtt14mIYd6YjYlO1FZsrE0uWx
u88Lq/haeRweS8/dUiYoTXaxEB8WG5DwDjoNWXsV4LJ8VUiOcy5xTGwU7u1p/C2V
ut/s34wK9BilRTY0Q95W7d9HIuek2EKA4/ZwltTXv3xRWXt9HYlj1oOs+Zz6cAk5
ymJJL5FMs+B//y6y3eIuYL50AaK10TSVokqMQxaDxf4pPDGHieN1s4X6u29Hjorh
kgxJfwt70MYjuICYm3PVtHu3gKsdflfEabcZRMI5TBnKmDQDlorOB7qPdeWLhjE+
/gH2c0I525kbjozluoasjm8YhP9nW6CY/RK9r9F/wnXXcOdzVWY6iT2rkiq8ybuD
z9JLybY83AM26iMevjjvshXzlAAHCBQ/1cLyI5iH0GRtLBlYIAcZ4c37pdvLRDVA
8HmfFRTStV2TsfUb/jezHSXQAYuVJZLwLPTGmOwrB/eqOBlXJngv3bkBGpcU9VzC
64MKj3IRvC2EP/7cBhrY4PFlXStqSwo13fgRH066WS9oUcYVDeHxN8/ANmkfOLTV
NoRc6N2sVENsA+fma89E/2ZFYH7mmH5mCtBZMCFBs4FQSwCJ3vtW3rj8Twll1qHX
mgckf2Wi/OoDpfZWwyPYFby6eqnBbAy04q7nb7ll95fyhFH65dLJhOYGD2VKEyEL
bEcrGYCoBEuI3qA9pp/GZe8In6+JXOF4WcePzFYimgOXXLvtThBibGV7nLApysFh
RA7nMoHGwrgzs29FADtwYZmsbMQpvPuKzR17I0HkK2Cs7M2i2ClYChVrifPoDAn2
bhy3CXxZhnWnG2QT5Ond3T0M5tWdVIze+JJoaY8LaaB3e9h0CB8MHHc4QEAHmomJ
sDDKJnGNPpDZ8XHl+vGMP83zqKH6MqNQ09p6qLISJZbhlG8U2b77Dr/3nxOEBNXL
POjQRYfp7odUnJzOPEHx/6XSsSLicudm/Hyo1toGUC7AXKvnuj0s7qDf078AL+L3
7T/5S/cA445Cft9iGxTnkK7VGKst0cgtfRJYAr7nC0+AvlhjJ0CvEezxCAgJqwqG
Tffd7Z/3RzHFpclVMNqM1EMOGRp4aHByInfTl4SUTGF5Ipm1no3L3m+KnlNEsFOt
t5qoCojBEciU4nvjNUEQdzx1ln/b5iUk39OswTPejZ09I3ctSW/lc9oIFTmkAfGW
j1mWBfACS6N0rQAyCLF8jdD3S8t7JoNAoelwN2NDgaLmm7Htzx7weUyQ2Wb8cQgd
7Vsgdz7vFCSrZeBNQ2tCWBcRV1j2C6wcakdGNIAR6iRua3oyCNmFQPDmFAbyXqiP
ONm5YwP109rM++GxN3ZnsruKwlA5e1Oq2KXUNBFbXBdwc5Ie48xcJrZZdGlN6KbC
HN40BpAQ2uv2wJH0aErMrRLQ54sITkT25Gf1lTmDi/oiZ7T4BemV9/SXsU1nTnX2
SqC7+7zpxEkgUTZjgOVDbLxCgrq8nc0BuFJdC751sv8r1scmVIYPZZ6qgPn1dL1w
Y1U6IPSvvxQWHAn7haRBDnV2nABaVX3z0d4loU0vC9caCKZ68kK5P//+ZrKeUZ8e
i389rgyfCYSRa+gsSQgbICDifWWHFx2UUXnXhd/bvt9Qu1bP4ZZl47KIzqxZASjD
+sYVy6sxHhZhxqsAzSuSwoEbKXETji+E/Jnaw1oW8Za1EWopZxeZE/e/kuvVEp+p
Pw4KBTNpWDFLD0b0+TpJQNgxxXfjnw2ID85i43QLdBSGQWHY2WRvsckw0NaPJhlz
3ThPr9lOFOfM64ZGBw1BtNUg+FSBXAuEWfZnkQ5If7+g2bC7ymyuUVQ6a2ORJLoa
zUT9t/1nAt3yUsDuCXonA8d4aMJzVOLFXfKVZG6dEgBGE/KPicO6FYivDzMK9CiY
o9G62LBh7i4xuncEceWgCOM5jP1/u4PBLIynOUTAbYR/X5lZrMQEYvaFKh+uz+wB
WT+Vdyvec8Ko+Lu5VVh/yLySL6chrTS/Yzg5ZlWf2Qm2ICRPaz2GyYM42AqpIR9W
eZBvjmfsSuJPXFOBLJAUuzNYJJnxhvSoIk47YGr11omMyyyRhDUoArH6Bts00XGy
CT8FNWvyjkkeVi5D28qLcv6ACCWFI7ZWmfdJQm0h3Un1jqYgMt+QNu257HS/xz8h
0V3F4bZlOvy8TJw6MgvOiltJeerljSZQLGfAGOcQmuX+59szsoqg7KkHaJyduU4r
mMLyBTzyz/fZkI7PVazvUwRTmCZYWIOSB5yA7dvf4pse/DF69fqFYv8mC4QaEdBn
EhOiKsCiM1KgG6Z1XmpC+xJXyl/DXVkdtn0TTps+jvAsqr61z9fTraCluYzU9bUJ
6tO0ITM88EccD3CqIAIsPT7fSqg+m0/z6Jx4r/mGKoWR3lipq9UszQiBiKdL65vu
RNrwRULzp2qnyyvlOlI3gIt3Gii69VdOoHJdIqhtTvzuZu/DwWYkP5RNZJVGSO8N
8XGUQFVQfBmMc/oTjN9eeeInKgDV3318VlTrJu2u7oQnYuyvnsyD348TlIzJS48t
t4d2ertvdyJtW5t6whJuZs2fB38C1Fufs3u+wEJpSitxPNXPTtGdY+mnVnWpd1x3
YrX7zZJOg3wNURmmzsEBEM476MZ6EZhxwrkJ7quFChFbBIc/w4F8W4UOA8dU5qo4
W9SNhQ+1DydAwXcDq5WsZh0VcQcrHYwiSOfiTyTY5oMtkFVKmK0u6veBQ4NbmXmH
YjoJlomidYOGt1Up3gD/N6zEp+tn227ZusfMXEsqfFvAr9m7vTh2euMI37VhO/1n
jlcwjt/LEFmsPl6nQgS+X9tDFSKj5Qh6Nc+TORgf++sIec62KM28VgCwlI8OkHqc
gD3PBDfQYGMC321SudK0i38eGEdw+04RGH2lIaJSjHJ28shqknc6XGU+vsPhKrzm
87bP7CA9VNq7kVoaUcO2Rl1G9laOFplQSlCVfkdt4Q0KzPz2fdtt0XKHu8nSK4Cg
dZWJjY+evNrnmHXAx8KrYLIBcARbVKvVKuPd9kQo4q4Xz/C3oUFKkb7GvdIz0nBF
8ZwUDI+BFjyqdhIEH81H+gn+X7A8O3zV5je4IB9Rryb6yDxHC/9hviIDVSuuTiHX
/3f/s4EiqPfmx9IlNmVGPPdtZrwIsu3x97hlnq72wL/IESJET8/uQw3ythk6T1zg
wUZAjQxgL8fUrCJT8AexewrxDk379GN+oYemaXKtVLybjp2IfzZ5bYs1+9nomx25
yuTdefEMzCuXxeIOkH++zUwZfiE4skX4llS1OMVh2GLpILBKu/LXCZ+gfmyrf686
R2JoHIJ/fw4VRwpgPhQ1brfUMeqOlWqaGBoMRpGg7qqyTLiYleKpR7xKchQM87bd
kbuswg8GFMvaQ9Zz1j/SgE7rxgVB5Cf23vIfoJS+BLiZEORqB+cNE5ugp+qDS5ro
c5zC0np/xpbmNXN9GmHpLbZ3LePgv1dTKwgDPiCb7i03Ka99L0DVauHHC4QbDsVc
mLyWLR8EP/Vdpr+bZMENwCZKOSblcARrUEWZ3BPFVkHn7SD+d22+Z7Rhk4ZCrN3Z
hjCjoz0REv8RBOOrO9Pseyr7+Mpn7QkfalGE9PADcnJwFfRZ/KB3CpF9P7jV7le/
AmpEVfdsJuTiKu36sH0qt3+Apn++l/p6zn9DybP9GAGO/NOJzbcQyLy53gl+ahjp
/lD3B7wHwcub+Bt5QXsQvbMqXpK2Te99Ofx8xEgQ8VEufwx7wrdsi7Zsj5lJTHOp
bPAeeUmcZPvQx/MbRq9BNH6RabarbA5JRXLvsFi/QXj+Gn1F2eucPO0FuXEXKoPU
t1pA9R5iyiOYsqhTE9gzSJt86potne5dg314j/maC1RI9deaCimCZBhk4KZI4AVs
a1I4D5n4ebyQAIf4tDN7GJVwvSgY+Zv4wcV8GeXdMYN8RuuU1nfQ1/w1t0wNFyYX
ElQqk7xgT4uf7rBiHwpYMdF+XP2hlqcgRR5JhH6ockALQNwJsF4uNn/+0GoVW2ok
IxdiRaXFHkgCQKbHRehmsFIvHcRmg9Q7S3tBM3Vd+Z0U7VcNEch87D/vpMdywkI6
iTLk7hz4Va2t0tlbr7ba33RT/VlpdXKrUr3mMo03kiLoZ3hBeR4v4g7yG+z4si0B
1qOOhR3B+BuSsyODC6Xae/4iRrwjirPNHyh+taNBtAjqVPvnX8FkyrvInVvG7aMn
LlM51dNIyRz6MFKiugeUHUlEEisjpm8A2VsDhULW+DzKf0epcDPrWOtBbxbZm6ue
jcqTqWt7veNkO9T8nkXKUw9+WD5KtpF5o4Jq1yCv/liO3n+EtFN6GAEiyBgyDkJn
krCsRxSwQ0FuvXspuKZUUb0ZtnZyPF2PyRh1w9SxS6FrdnMKyI03I8Qw8A/y31xs
7R9o61wuBoo42/nOwMLhYBRZlPlUXIjCQbNyUVpn/ZJmZibh496Fm1ZIZIW+UpUf
sTYW9s2+Lak+GKonXEPfxxQfkzmkem96XxuDKLeV2wjloBDuNTb93Y0/aQrSF67U
bRi7K/tGajhqlUhsNruTfqYbg/koaipkSNeR40//nLdXA06rQrtB6mbCgCvw4kHR
wENfUZdLAM1+OlpSxzeO0pV9nuc2NpgsWrH/SSuot9MGW6iJ7/tICa2K1clPHyPv
7J9kMOCWZbIB+1O7B68/f2Nldc8+B8mi7gySJ8vCDlukd7+ZI7gpUXE3BCVra934
bXg6eKiacR75QScCQSM4e4aW9e8xFIOXMzL7b8Ax+oQevMV/r8M4ikV0CerRltdS
56tPQ6vrqlmxUSJCjP77a3CZ1PfEb+EkhlVIMdy72f003DS0yFLvOupfGjLLKsPw
I3qTvVCL59yoFPa0mrEUCUcAnxb/rVI9KeOTV/m2K2b/7cOUdLa9YN2IXVCpa67M
K22NINVwwUXi0A6dbnomCUxra45TZvQx0J1x0pjpwM4w1vflIwLnlDFQxgvahfuD
yVZOqL2CS0hKnyN5bdF6V3BXgcs/tl3Y301Al7l8Hz1Qt6ZBi6+0dPOq2futEvw9
5SFRpp9uhIa6dhc4C6ztTy9JLVG9TNVjCZk5q/4yio3YkkFBwAHJwzBndnysPQ5o
f3hM70HiuopY8lLiK4KxAJEjgx9q4nU8EbR6GHgYImNhJDTX2kyTlLmmx2Ak1Fig
AxhKxD5LIzjECcOB13avG5a3yNwmBF43t/ELd5hHLUyRWLYCSh8lVUNXN0nmtYhi
lLLjL1y2tE4eVsiL+dpAyhEwr5zq4mXyPtTkrMeApOSEGeWpc1u/GvgzWZ9ihRRU
M0oO3DIe++a9nyPONiw+NDAGhCRwiWwAbXeuVEuA4jrhB1s5OB8PBUsGHj2iTmtX
w9zEFY6/nD9WJVcYoCbz4suK+4bwbFMbO29iJU642neE92pborYiOVk5lh1uYEkk
XlJOZOjBsvt3lP2E17c645QAV4a54dbvHQ0dIhtticZQ7YlwRgnzJtpQXG4H6MAd
zKAnI/DsDe2guTtfLes76PagfU23iN6TmWW9HETIa5c4Y+r2yJdtL56StBE1lu6R
LIJMOP+9RSxjUp1Wu8yotosRewa4XuOyFA8fPnos3JlEZCvT0RX+HfvKGoVpT0OT
Uhhv3YEhzZjxu4znte5GSCNaZDTr02p0VzUIsPdYlfiCq9W/FF0bg7McSuv6GjCc
9DW0cJ4NIeBZvWNYR8i7DPNbTFbYVvyAtl+N3t4pIjW+pVLoh3cxMmaTvUPnl/Db
370HGc0+Mfw54hr86aDdNhkB/ZEOPH/9pecBdeWfTNYZ6y+JYtzcD3QIRCA9vWWe
yvGFoh7AIB3MbTQFyIN8ZlxuDsNiyHUZyXSUS9Q8I6IAS5wtODK4fz6fRnDSPzcM
ZwWvVOOtmhqXcRnbEGnccAyhdBt1IrPYr+bzxb7hFAI7FbJIBql2j+bgv42b+Jtf
QZqdD7W8Q5F7AGJ0AI8/o2sfbxACBQhZhGkUQNubTfO9lgEbtxToe8CFI4JUbevA
jQO+QCPEbXhpYgUkC7BKFSpbE3Vx0aED0mhlybc5L8xI7/z/GzZKq1ADzW4qV0RZ
C+a1rMR2oqLmop57PZCoP9D7pxPOBdHQQFN3EmWWEItwvccqzSHlJnPYExyfQPO4
aDaBN+0hNg96J+tRVJs0R+0s2Zk6XZmEn+m28DdF2cz5eE+lV9orr/mlcNaxC4iC
TkVhrFHqYU/2jsqaqsntqnDeluh3tkX410ul2MAQwXO3FeqUVfNcJY9wsJabfn/d
iARtYK9oqorqQnfh7LcTomv0bYUfy3PV7BF0bllYjyn0jGHyG5pusexcsfoOnxR6
wysA0FCtoiyb3kjjQx5onn/ivZ8Dm7gLDXnJMlpdTU3d+TKU0hES5L8qeRvZ8SAj
xjAeQXWhs0PSdeXJK3LlRH5aB5jlZcpu2pqYWiFG0k+3dJ4Z8yh8o5pgkQvFaLMk
JExqstU5qzM+mM7mvx3PMg==
`pragma protect end_protected
