`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dRgFO4NYTPppPKD395qMz57u/deoELwAIF8AA4qHs7AW6FScGULlxWNc2CINzTq8
pneEgwpJi6LJGBkAT0AJ3Fkuz2+FhhiZA2lOBSOurp2jTN/PRIE3G2pqx/QjlQlI
ofv2AB+q4xCPWlIYJ4relUay1uyfeh/WF9k4RVKvalY5SO5v5lNZ6fvtd9Wepysb
pjeI2lGAqo2RKVPOqMyQsmU6+kaErCefheg/eqUwvqPvTxM70buucKBnYqWt6P3i
y/p12On5wTaHk8P9Nk65FvuDcajgeymncJC31oK8paKq0f4eB/lAFAHeMggfVtF+
rTZZJ0UGCP1KGeeWXWGz1A==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3024 )
`pragma protect data_block
1OOUzBFuJ0AWil2rYWFPuiV3OPWIDIxJ/Cs+7RsjwW4mTNW2OgfcQPd8e/fNLAv0
qW3lIt247xzS7LXTPKZiimN2Ohg2g4m7FNAHo45lBQo9H1+emGr4EHkALHY2U0D6
jmn5cod/+Uz0MN/Eqj4RdbdNjZ2/XNRpcREp8BV7vCLqPmZ0ZRTWHfvHgRiVXt7o
5NuCwPjumED6q1eL3msShkrpF57r7vqdJNRai3XRtlnW+dqndJY2S9NmCz69X8HU
gfArP77Sjr9NlHXdPFPRdCNYjMYMzYH24SSvqWDvQgIOZ6OjoFQ+5RJTXp209jd1
Z5Q7stwNUgfyn6NW5PbwT+pWwL7l/8mtgP3nchQsqLPujJUc61iBga5ZbLLYnTzf
i20MMYVxnpjyF9crS6lpdqs/6mrir69X9CqI//BwseUk/jFT2HWhfDO2+GnrkWAO
Fw7WLyNMVEffJRd7MbQ6nbveYk4ekbRQ98QDvVFNMVs2rMcikFNSjQaHgGVGEqqq
VWWC9TnL1WCuQOrwl4IRgU+TREh4j8ieh2gFoYJvdOHObxgBGSsSlrGoTTVoq932
fhkTKq718Oz7RBNkUcUF293fuf5HTnbQQcQ4yb+TrW4/5gZA/wSeBICl+m2Tp+hO
dIMobhcpfGKzRWviEjvysZ1u8S/Ff/zim8T0zA5aolfvWhKLP2Jc43I80VulQNoh
YmEkRHHHRWlNtlYX6niyYYDnQ1NfK8hRBAshLfox8eRElh7GZbeH2pS0h4m3yySu
JkV1HxV9UWoLPta6Dey+TmsalidntYeXjMNZHm/XSJp43/PRxEPSl+ww/cDfJsA4
D1Myv/ljTbR2UzbfAeTY/XxM5lNy+/84MCFBQoKibMlMJ+DvVb5fGiIxbhpsnsDb
APxht2n8qFb/844yAPztDEx2KKX4LEm5EGYKOSUFnGvzSj5uck8LTKPsC1TVMfHb
xRzek6E0Ct9pKguGhC7z6FuLxysmja8seH+oDwAoIo0vHDnSnJwvEStULG76D4QC
qnXociex43w/T7n1+Y4njEcExplSbA1rTP997nAXQpSdPvp6m6caxBqKUMO6FwpN
b4MroTABxgxVNPjY2gwNf5ZArJMOrU1U1bOnI2ZSDpTx9xRRmn65YkVk1Rxkome4
Aypzev7FOHMbbqEXwlQ0Xx1YJ62Ib/fabp0SPlDi4JwQFIRu7GNUzYB5jMdm8U+7
jwNiyo07yH7ZlcifQf8sVMuFSChG/2e53x6xv5kxwcNrJ3z0FSduUqqRX48G1JkQ
qvq4pASRvD000nz0jyQBiGE4whdvPV47keMZQR0ZyOv2I1ieEf7Pjwg0PIM0Fg02
yAFNpRRjosgjBWy+04+LzYtg4Eh2FGfZfOG1YMWmUvisiFgFAhU+dxFKCOsdd6TO
gnLiWwBjjSNf2nhE6lu0HKNkjNjFhwdFCjRcfc1oLybIq+Cs7TVCM3R58MIRvIQ5
0fY8cvBS1JJX0bdMW9v8OTEbbPgss/oJwrMx4X8XiYVoo07aj/wc83w+c+u1eDRS
aCKlZAxtzdg9m/uPm+wUbBjS949/AeDiDCvCXRDSqy8AHAOM5knBa04RIUBXVzim
afyJWT4hHRgqZoRwJfkQLdyaXi7x/0d9BIUOwmT/EzAfv/a1253VIqmblkujAIum
qFBjv8SHLVjFbgk6DvCUV3h0G4VrlkpVjRrxMO70pAiFI3OD1uTfnE9HvA5pq0eh
Dq9CH1UR4W9f/i1YZajUDWkHmlax+mCrfMDgq3MJDSKW8ZpN9swG6F3IitotiKCE
Jzqk0K/a5DT+8F7bcCfYNS+dfgRtHcQXy4W18NpSZEN/HsA5OoYesd6GTo2QECpk
1b7me9/REVIxzL/G19rA5+UUdzc2S2Fg+ieQjJLyHlKutHNIJW7kirskqzrX/bJp
+rFBjGsjE//5qg8be8JcRlaeNeEQX6dYg8IQPqU/yl2Hh1SsDBs/+pRB+kDMisTq
LVH/vGEsQa2qbWOQsOnTTq1elma4iGxofi9R29GmMjEjcUE43sYUD5KZ40AsluZk
qlsUqJ6vOqTOn21C5PJp/IT0BsOMLq8y7N5XcBUjR2OJMb7fy/WZy9tP7nT2b3dM
1Lahd4WU3lG3252lHghRBhfNUCEWWuq+Mrky7VcuiEuABpof2o/dGsMSMdyvFJ+l
BvituukXYDihtRKOy3fAukfkqX7nc8e9aCEAyXSfTjkN7OjIBSzMXQCuM+tmU21k
bIkcxWbAMAjg0yURYtUL+yr7tLXsQoK2oMEq5uDYZN/8LBx93Y3D2YDetPcB/enn
oK0cEfhJND/V2BQZ0MKyjLFaxE5GFniRFCIbMIc9PHQdEg0UmQy5VqRSCNRz9QW5
l+CTcwi1RzOmup69L42RnvhEQjFv2Rn7KwO8yNubs6XwUJvD06Wnw84waSC7iSJ5
wgYEBR895vd12qZ9+h4rGcHt6HGtR2nddgPCo7aWFAFF4qvKpXWZTW0DDxSIux9i
CaWTmxXqhE/WR2J5j3iarBqUYRQafC4ZslAESX72vFvOLCeXhG8mN3GlxjGlHuJV
gsjFyoTmkSoxmxF1leFK0x8f0Ig7+7Rr7r1WV+u7qwLSYPIt2ydOfATZ5JVds/Xo
jFO0aMulXfU21rW5izgok1cUgYmLR5zi8N3EYzYvKazUjaRBxhSb/NO5USF9ZVU1
U0fRP31GNUOogU9TgT4P2yUyWvMjp7d59VWx3zm9mGzJubxIdrCMnfx+PU/CNy5c
pa+U74+RTuMl+T/Tw+XMv40uu7kDnSuMqVBMPVqohFrhL50yQ9ckve7PJy029dtB
IIkBPwrQWpqr+BvtdCOFmo4VmnslZVwGxl1nn8QKGIuVUNvn6fhSK9AscmcJ87/g
i0Pex/GcMzVBShHCXgUZwO0DrmfSmfAVdgoOUsAGNxV//+gZ2sOmjHQgfj8WxKE0
1kA1BMXH+mFjlvmPS3rS1x1bh3ZeJ6EMf9A7fdVYWBbM/WJfWBqXCUzahwISj4uq
sZ/JDAeQwBQisK9Ov6QWGXrBRVf4Qm5zFnnKhHNktcAxRl07p7awnhqzV/IKy1q8
6yZHJ5m1J/RTV7QKVIAFPLJ2U+UhWS/MUm4f1+4K7B1nnCC4OUfeSabnTPghShdB
sHmwn8b7f24jjJ7UdZSW1XZItPPC06u80IAC7+2Tr1BoR4t5x1Ykj6apblpTDFm6
bYGhCGALoPYADlPamSFv02sa+nPCNiX81/I18ulMu21pgO9/cBimTnNs6lLyiZz4
cgdn0DUsaq1/ciO/t/T7j4mXBuxkOKd8vE5wFQZIOGDEqvBpNGJ23N/3NUGyUAvO
kbGuG4ZWS53wmasMhnw6YzK2uEKNZrl3p/luRWdNfakX1DRNyTF226q7MAIf2UFb
M9OcMEZKue23/yAwRVrw+4RuoksAaCQrgy8R7McLYhPT1L3TKjDr/roKZQkVSX51
0DzWV4kABsH8sR07bmF5e9lUygDL/hFoUnCuht8cT0DTKNfLu9Rcj37HCYWsHyd6
cIIYwYRLUWlZPDySka44z9/RpA7SYtiqhVFLbn1zlAkM4JqxfQG3TXv/mBHXIiqd
FQrsmfDWPcMCln+EsWQcmdHTi2l1W6fI0eW+Iy441EnQgXuuESFoVzurCb4N72K6
ZkhwedJtNHrmEkAxMCmP5f/pMfRM4sCRnUEZ2hv21t8BcGnsw37/2AF1XXUE/4c7
5+Vn4b2VFl7AeBlCtkjUWah/SI8rBjUDLlr/F44zLevSQ3Ht3R8Vm5JIV6/3TW3D
XuBIefhrVR86G6VsiJF7qhTWGWKEZlxjkdaGesXXblDqeR5Vj3i/wTn73qJVkywS
Y2sXx8kAfOmXx4GmKXqJFoSQB5xEvHiH91k50YeRpXboQLaVbxhusplB1hSdxFtZ
i330X2FQFfvEULA41B8uuMjS19cgbGjpUUdcISiexwylNkecmEJDZoUvd9Id4A7u
oDVMGwsZo8ATB7SLi8pn7EbAWsAywHgulF5CqL8StkI+lT6M/2hcaa4fkFFqtlGy
`pragma protect end_protected
