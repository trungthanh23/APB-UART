`include "apb_uart_change_bit_num_test.sv"
`include "apb_uart_change_stop_bit_num_test.sv"
`include "apb_uart_standard_test.sv"
// `include "apb_uart_strb_test.sv"
