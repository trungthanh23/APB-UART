`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cK41Ime4nu8UANlJKIUUNCTWeQi/Irhp6nin6pk+9MxG1y9sU8KGqoNsiapoI6F8
Q2jSGdzgG5zVx1lE7Re+rD9jdqXQIcBeQLMCvrHbFLsWkoo3CNvcom0JcH7RW1mw
iItWO02JStsIHfyj/Yx86GB6hPQLD6vqbCSmthniQBHMtCbZ93KsdlM+kmVwCKAt
pH6ccDLGQXVORAoFBH9xpw+hVHztF2DErDXAHLakt86Tkwl0j55x4DUnrbWK+naH
qWKzkcmUobxMkgIigl6qC8WTl+kztMbuu/yVS2AoDOJdUqTHQLU6motUot/i3R5R
+Ey57Rk1LLtX7gfUYXZuAQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 352 )
`pragma protect data_block
MuPDDRVgKWj1b4cW+C7rS2lJS/i2ecowSaiRNoG+qd6MYH74+byEtVhX3+lBp/AP
o3MgoWHea3PHMlT8owEZnLk97F38ldMvKCQpdSgY8G/103K+O9vhk/oV0PEB3gB4
KXAWgodqRwdvuL4AUMl/vok+orDyAQyJf9+HA4TgY+maAv6OmhjN1XZtJ66t5p2F
GKqPu5X2P17OYvNcNdV5ki9crI5Yu+5RWJZ1ebNsfhmoq8Ew21E0fVzP+KzFEL97
9Z8KbTdIhXyRRJIBkkkvWHtyEAnbILmNyIBtZw/Zz3GpwwxLfxHzdFGW49+7BzaG
kdaw7N4AcfdeTCHUqaviQgoieaY8qCSWCrsP9s15uL6hifWlkH18TDpxJHSzwEnS
iZzRN2eIDy3L6wGkaK86mSCz8xKOIyxqdXYd407R6s+nqYuCzRP2zBczjguK9NKk
JBQLk/0I95SnbLDaBqd4yQ==
`pragma protect end_protected
