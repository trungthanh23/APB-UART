`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UbZVIdTVfpff8WhEvK3uNg5s6Xvqez87xHxGKkvQqxOtGT+Ko33JaZ6N8hsqDYm4
rZJltmg0hHVfEVVqwmCXN8+v2T3LoSl0dYgSDeY+yKmQlkcDgkKrWXR2ZFWspouD
Sx22lDJ64PYEbmmWC55SC7ueiHE20O9+HJgEe0rLCUxl3XjW3Io02FF+8aIs1Aky
NZtyEsX0Rb4B1u9vX6opr7a54KCVCPC+AaUunKtUsU4r5sIHo7igXlRJl5vS1D7T
XjPJvUWik1TJc6S79/WyoH2tGQQE6ZVItQM95Qsxf2JZX2ruqpbcmGgTDz4t1mFN
XXkM88F1x9lmWXZa9YUzCg==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1744 )
`pragma protect data_block
oTX6ispHQQAFzxGG3I7b2dAseAK6pg0JdqQQXUGevglAxT47UehWgrlLtcPIwhoW
Doz+RiLW5z7Qm6zMLWj10M3oN5yHXHQZfb1EljO0e7b1ZbqEtY0/uKuVerVL/K3f
JHz09Xx55o0WAqBlFYYTD5g/Z2dQEK3B9cJyJjsSk3I23XlFQRM0gkcHhKmlVuhu
BjHbr8LMxPN6d7i0iqGDs0lJoOpuEZWPc1HbknJ1yu6Re7O5tcrjhzJuxLKQrP0m
xE4PoZnX3/kgfXxDtj1v2amfIbF2SAOfkc6kjr0A/b7Dpnzgw5tI4/BJPeYWSauW
vXYKSD32KaB7uCKZOFYIW6TnAm4sPiKyrGANKuwNdQCkKFnmyIm3QAx1Gh0FNnVO
8oCzA1TvKMw9Ve/ZaU7ykf9CwefJhH1BYjbKFQPOoJY4v0fCGvC1tROCzHpsBvNA
JcPF9uOVerjbrXzctM3v+K17Yp9ooyVShqMwd4bKDpMsFnH/sPXSosmSf2SGqxc2
s3DREPiqAEKQFS7MovZvPs/WvsgVvJHWww+CGVCK+i84262J41dgtCKgY29PAnfd
aleFpV8/yO6dZl+tt7qn+JodLRMawyq1rMAMl2V4L1fYJgVyAf1zN1maaEQHxMXF
/wFCOsHyP6KC/2TiUf5SM+pLRG7+8a1DAqRh4Zx6BCsKPG8B6XIeT1olkmFRGkcN
CT9CWx7rlfgNup6tviPdV8xd4QGS4vZ15PSqoNmlbTVjb5kS/cRQv4BkY2KUvyTX
zBcqCeiiuvmR0gz+bhzcLHjTNQIXZ3fvpShJvOpeo7O9cB/a/8PzhwiR6sg3Q4zv
PIlkmDAKKBGRly8wYuB5qycCVc9IkOwfkYaLEvCOxv+YYL5OKreQSSJbCFxvkyzj
Jz8xk9FvfeUrmQOGeezkRZ7CNAFTjgj0l4SWOGdCVdjlgK3o4VdJmz3urfLuI/3I
ClSrruHUQZq40Ps0pv39EQ08ZSmt2DagezXRGZLKPQqcCAw92ybJT4SjphqMUV9C
93bVANQSJfJKrySWNu5G2DUEFIv8EsNKgL7+V/z8crVLUxMLSzllbbQWnlc3jXKz
fGFsxzJw6qZZkgJOm8PnHRatM8/RxDa+Yul8hdWohuzPskoYFWWR0RaWiGCbY3bq
q1TnTtMCWgc/oTaj0dcC1L+e9S+g7RxVYotllhWob1MIiwutMTO4yHlIL4rrRWbM
C/KS85LSPMKZTpGgHkjxrTh41/j/QIkaqjTWDMCquoOwqt9olBUZiD8kexG45MaZ
2qss/RhdOyprt7DVSzIYIfbC8zscLQiiWRqudJ8QEBpOhm98eLh5HigMirWIrfm1
zKZA6IBL+U1Iom2UWQpuXqN9Ry6oUFhe34duOLXpEbUiqPOUDCD7a9q31beRkPV4
5qEz1lV4IcJWe/BXY+2839e8cBFIBTrJ2tYX/xoQ80gOVnxHUt9uFb9AHaD16Vqj
5biUQ2EEg8J4qFATWtbSHe2IGo6//NpV26b3Mx/QIy3q+t12bYK1b2BELm/ov/c1
tHdLTzWLH8tF3rjPDmOBeIR6g5yxxcJUgcyj9Iwxo6Nvqpk3D194hRg/T4B8Radt
dZAKKbyRLT8rYbpSLwfpVRPe+0s9en1udbapTquuOfijKHPL5+ZCObQ/JXkeuaiP
hUnijFV4uXARcMDYmQ9H02/pUu70xY33qXNhHxG4drbuJTAzf8MDShDa1q4Qkj27
GHZ31c7FCYtsAtxNnyjpQpt8ge/PSsxD3IKw1UI/47D3Idr/LpIFmwchou27Suku
OdstXnegD1MRmpudBzgKlIm5cWTj8I3gNs3WOLl0DAsDKDlFmdajPbTYr1u7jTe+
vqjP/9bQDFAxK3nXC00toOaCgUsEY4PT7k0kkdvoEdeeheRHaO3drjIPwoRXrfDj
umdPfuecIQJwxTxhuB57YqNNA94qTM66+gWm82DjJOy/TPoEHbxbLu7OUfqvVB2J
lkUo9g9rivncDItQS3iOCvIdZnyNdEuzcy/NI3DqAoKCu34OqBy2NBZoPOncS/5s
6sbxB912UZ5DbSTXJ0KXT44wj9L4eQqJHHx3svIonxHUzXygOYVjcMHLfRL+2YwK
vTGLWWSpvlOxZf9xAMocTP3E8rrNlHpJZ142LNC0N0AKSVnRP39kosCqCbCgODK5
SkD6+jnEaHhZ74qY9SMH7cBHg9yRKoVtCo1h9rDVjsn0LGoFcQPzrpSruClY//Ms
LGYhkq9IO9ERiRAXogqXuHjuEQLwa/ecVPvNtU/3xHC4ECQnXzsMO8mZDaZz1ElU
hgHFTOTQcOZth3SPXusG3w==
`pragma protect end_protected
