`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
F74CIb9xIZSPvH0i82yzFivFQS7kqGyQcjlnbAxQ6pTTNjJ14AOo0wr1wUAOwX6R
ULXjW6n/pYMSkkqNFw+gbGiuEAQSswD+kwCUmf2hsI/VIDIMKrPGZkZSpWssBp2e
wECi8dW0PIkPa/l8zfZJLVt5nnVKa2gHLC+zraiHK+pq5MN2Gl7g6R7z81LeiGF6
16QUB2kmGIMJmSOQvfXWFaC7deUM1Iie6YEDmLi/+vvLXzsFH0uWJhGHiKsQtcHP
hMAPFr/HlGmi5XEa/ABKYRTJ0axL1V7Pl9mTU+XjcB611QTV1b5k9X3uC+plw6+9
ePVl64U453kQKXhLBttlOg==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2272 )
`pragma protect data_block
j5mw/1kYOcpEaxdx9bGwGhY+KkUIDBHVQukx25ORmS73KTQCw36A9n00N/4kAJ5D
WxgWXRRczox6DMYY3vc6rs88YhCOtas+BfZpTwbgYwaJFl0yRbmHxxIO7ESx/gIP
mgAVESZJw/hwGA1ubyAztusSdZ3S1R83yC5vH9EqcDwzuk+y6vVb31bYaitcNBE/
b+G1dcU9UQ9PCD0XsDIhYFTLmzOe7z3Z3yz+JDIrBRqlbGwPFWQF1EnlmWbO9+mT
3TE+f8VqYjg9hCQpCMgCiEZi7Asu543tdDojbk/GJWpIQQSGHOdvHO616MWg6RAT
AlQUYNZ6dodSXZdnlITxn5u4R4nVVMB1dnd7ogkpMv9pr1CMsVEP13fzI9ACUG7Q
KaetBF+mP7RVsxVGDa6EiDr56c9bkT7OIaR/e/vbi83IZ65rTDm6Ml9b36aOi3/R
LqLVHWQrSX2Ygkh+MAZWJOaLdm7iKOW3fQxhSFGtzoe0W9FWU7O21rkEq8SaI+p2
TtOLDBw7XGQaVmaRXgh3D1DgG2nGnzNC68FEK+o1/i7ByVKfzxbe87IShoosdTZ0
QxtUxha81k5fX2cwarvWy8Yd+DlQeNxN2hgWSXMzV5CHrLwu0cArlz+cSGMA0qYF
VBPBcCXYl5UzQ+QFmJJteGy3O2m+u4EvznsiBS7r4a5XjqHNXylF5nw2gWN7D/No
GbhsL9k5KfjtbXXMAwftEltAN9WrRhWliAGK8h0FiWtOJ3d5Jue387oSSzzCIWBH
QHTpt1u5OqyS0pYya5aS5GAdfxVupQuhy60NiSkGYxtHYna45tyAloqimSZbMgYr
7VjiRW8bLeLhfc1zot60unBTZZcEMuE7+FbhlS/TnBy1Pyw3lS+GPwB+D9l+CvJU
SC/SfSz93R53rjaFGxt8cOMGY1783GBF3YO8lOFik5kvJfdEZBPnyz4BdmZuw1Xf
WjzczRrEsH2/Mvs3CA0rGFYb5Ke26Laa2pSM4dv2oH+ZQBe3yyixgS65gAGN2Xg3
yQK8/Mmv2RC/1zD6Kf89XjXOcTBcAKcnT7b/QUk88poa+PCGQuaopQKJPLo2hrf+
y0R3SenTTbw7E/yxKCwh2qrF+7U2ouoZSTzQ3ZaqNU8LbG4AbfE0zmeAVZb5Q/+N
aBjTzNaLshRm6wNFpmbpZfUUwfYn8lwSFlyi5/MOWOW7HwHd60sFUyBr6eFl+gI0
b6jWCCfmV7qZ4MbcX7QfYQiCECgZ9J0SrGzO3qOpjPPsxZZj02bexhMc3KEgFjkD
TaeLhFWcHq62RjiIs8JZXtPiOredFHbvgTDgl4QvwBNE9m5f/E+88aTOCThuM/vB
DHvQYQDjswh/79wtu9rN9bQORiLufB69MR23vLl3RTDtVvLq9uQKrWyk89j3bAHr
Ox25cQn9azanILc6/WcUMVNDYUknU6y+6nwH1XiBqacrdcOfdFf/SCXbevAlD6in
40+IBdPVY5+dQEYYXrOhPRaBRl9IFbLrg3OF3IPZlogC+/xrf58ev+RtffnDvON6
d/gUJ5u0TrUjE5yGIja6Bk4rfufFsia8g7bZlcL62Py3Qz9oIQjx9UfvfEtMGwUR
oXo0vxVZbj+FL+AnfB+yXbWiiOl32DAXBxJYa8c+usrOH+T6t3NK7bt2askJTh4M
/NN/m2izpDlL9wanScExLUpTG/kaZFFVRD4Oi02S3dAgrSminCnFdAq9HPqEwvXt
q5vBqkB1xhor+EGLTzijgkYV5o9od7EgLcpbjpwWPz89Pheyka118R7q9GmDp0Of
Tjgkfd14KMu9H0dOx3JzljFgbH7AKNF/LxWPiwjRjVXuwVqcCzSvyWxUWYYtY2Le
nfeNDEV+0w86jT3k0dOZ1tV4J24kyOBCrVExINGrXVby3pLpnB1riacoypAa7ReS
R1JYlmws7q2o/0mAnJxXGqFqRK9KQy+7LMTHBDaqAyEorg4H8sShS2+b26CARnUj
+zFp+MgNFg2aSr2m6HJS24QsOW6cesNcPx8VNRsc/hsEoLJtXHfAhyDOWHl2te8k
vis12p15NDXN6qmDGKMkOwmcq+LsFkLIKaLCg9PfzXmHR8ZvmokG/hk5REqAyIMx
Ip1AcM3CMZwL/aHeWhyloUj829UzMsFY/xm4MrGBuTVus72yOCdjjIYomycJ/g7A
s+rM1pQx9IuwK9jKUf7u+jBNGSamL0qqtVUDSAhfzmu/hG6xdr44FNMPn+JA2sN8
wkdR5Xlmn77qQnBYkmqR5PCLZEEW2URcgdslau9N9o8sVzZ+bgSoC0PH4EGuXO60
GrcAtpCoiW5GI1cAM3RYgLsdBEd6x5sptqMnFy3w2rBoxUWyuK8yrm717BGLzJxD
cTaPFmatMvlfs5KVLBJ6OONwzZtAXruQUKE9B+42uHODHIQIgeEwBGUPOh4rhBJP
K7z4koNgLtrnocKkpz8QUy8Ozgis28LUzMvo8inCoB7zzLum9YAbs03zvYPk1n2P
+hfbOpyHL/VhJjN7BSEretNFIgcBY043oLfRtSvmTHwBMIroKvJRWfoZUKHLWLj/
Zgs3lKm0QdeUf1jAzBH4dGodyuixEwVWNxvxOjETGmGGEZJwT9b+jeaS/edCOy7V
IUoozWZOQxCf8V1NuuiUIAoGpzVaE/+7XY3g70qmk92BiUMp1tHMraMOxRDacz5X
1htWBHxNiqi4X34dmsEopOs4DbzXZ9Fa/aYLa6cEupwDc+FyQs0TKlc40y3lNfOV
JsRuw/i3PYsxPYCGjI6vdQk0q97FM88iUZfloKq/hulbxP9df5/1ZWDjxo7YC5wQ
Uxs6X49xaeoV0P/enJyxVKAWjsYp/Jiy+BpQy8QgDpBotZ+fcs6whfGUhP06xU6u
uYoy4hydf0NMVG2tGlr3Cz5cofUBPzDok+Pmc5hNZhFers0o+mliMBeWLSaJrM99
m3+0MDt5HrC+IPIVezlGyRIWrcOaaBwmE7br316Uglcntpj5xdu10D20GFK7oWc+
tQAk9fg/iggY/zCqxrxCXQ==
`pragma protect end_protected
