`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NMeSZuK+UJcTR1V8Ch1q+xaJL/BJlwEhJ25gJH0v92qTzm0gB1DUf7Lhu+9CImAb
id/Dg+v7/pwQWr4keJcZjCV54K/ljHOs8F92680rLL4A5nEx+v2bt20ucMeGT4RX
3ZElLTacbRkIM8UfXkVc486LxPDtKcXftLxsyfdDsceNF67a2qh2d3KTNvuKIB0f
/99fd6EOLAhI83o80vFheXIcCbwHmy76lrKcANOgz1wbn0sm4Aw6q72IKvoZSGwr
9DFrJ8hSa+32lnKmI6+VgWikXaIz1+MVZxAUrH1OtXv8IbF36MWdXVwgwhlDQ5SC
E1yZZPpCv04tH4n/pYxCrA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2416 )
`pragma protect data_block
g3XjGse7rmourcMQ+b4pM8FWFgFU9XBW9VE1fqKXmP7cDJd+eVUwrkYtLrjPGPKJ
/bxfgKY5cGtemyZdPQ4e00CXXaYr1pnEUkRZDmvi9wOj37lq1gHcLYXosAhC3aZC
zs2VdQt/nu4uEyTp+zM8IbLkULVNWJUBRAkvg25c7jyLlSaGJU/nrYQZYoy95sEv
Ry+ygTIzshIzQ0AZK2uYldmaoq0yGSqutfZLIJyjB+Dch+s222w+Bd/g3HhGUw8o
IBKdyJbr2DAGFEmbbDGGi/53eLLoTCowyW4pD+LBNOI4yYUw/z4Ng8sBI8kq2Pip
SUH18q9BG8t9lUeHxmU0TFWZFgy7DojdteV6LQje4dgs2ZB4WuaeGdJ8+vUohKcp
JYlm0mAlSSaodgEtqQuyl9PpzhEHlyxx06Q/FJpHUkgr0sc3zoiX3WzAQXdXStZm
jLWJJIWeze14pb/cECiHQUp2V63qJ0gWS6L0MkCa89apx4DkIPEbbQA27Jl7ECt6
O/WZkOaQNh8WK84yEpsOcbE9ujyEMGPWZXSOUKEWOrXmQcfGcrV13kGrLIuvAhfK
49Nd8qFathhrQQSc2l87Y5jrkgGjLpl6qv7CAZjxzZtoCoARxn+lIm0Zr/uJePwu
kEvb/wg5N1flIPK9hR2HsdoR7eUZGSr7Zy5EpI9vJm/Bsh6jVcr6VEo4ufc+XH+B
iNZnz87h0nDfDo0I2Y+0Vvi9aC7gbOvC2RTzzJYqGQDGfDQigSePyRQuqm7pN95Q
VPn2trs5OYEXaLd0bAl/LN2K/WgCVLWMLDpC4TL/zgDtJJuuRkve9rC12qlQEx4b
mky5rlt5ipdUcL01gvEcyyMVJoV4pmpkMD8kAhJQb5zQxF0H4UGgghO7bMgC9wp8
nm+0Q2kdkhpctzFR1HT9tJHyBFYJnDWXl6IxkrutEDpnat42FiKRZRFeIcYCa/G5
5lCxmuJ/aWIHOgiyR4Zzu0nprpAyRr+jW4FaM37Yz+36H1oGuOeMyqMo5uH1WWBA
V9s91ryVoG1iAuiEMN6fXlKNQR0Q2H0epn6vz+n42eVnYmjMXbb7E+/N1N4OVe07
TPrnZFtZEYaY2dTr+XlvgTKK/XrOhUCsYdtHEBYTBHjIOHu0YOkyiXUCl++IFWie
sVyAFLOUbG6JfBJcEpJIDi9w/FkHb5TH+sxEUg2bV8k/80CtTAz8oyh6m3tTazWC
RTHI/ntN98fHKXlRJuItSbDGCY/rAOlek5L0/bJxoJ5F/43+9XSCSz8TCMEPCxl/
43yRaUfmhyOylb88sJMpq/FL4ml5aY4+dPFCeu3qjifXsf836Psc2amEwyPrLBIE
41oExze+dtQxBtioOy68cU5lHwq3/tQ4+odytDWZ/WZ0hYuNf0/cyK8rn63IdMmn
zxYKm/yP1qPk4VgCqIT83tXuwB5TOgP3BfT+q6SlF3PbTfRXyNx9LliRLvQ5Yw2v
Ttoh/6p2iAWZVjCxrq1HMSEKmCgLB4EvTVZ+j8UICMLw6zul0ClzIJUrgRJ79+Rb
DmQ7n5MN/ws31QKrw1kB5SigVVsN3eCe9GixDM/1FaIjA0IC21FJL2ewqI+CseaE
kcjJmjUnCUFapxHXhRa9Zxyt0VOFz9CE3KeWmWT1JidC+dPnZbrZZYtZ6puZWy/K
+Fz+ozM5jJ+c9Q2j0IsL+nUFV7N2IcrGYO9qRCnvNmSontpl4CoW+yFmjsmtAM50
ic22e49w2S24GeiB6dYN4DR+8PAjnqHkWeli21rJTN4EfhrX25zb+JgOygv6H+IY
CoJSg4zuWuiAKg0LFiipecyFcoJp6eZqRsaEWYi/1klaCQA3CpERejh+xbbgkWqf
HBSE3BG3qF096s7GexfmT7p58qzklJ6/maPlyNOvUB7NjxYcuaTLa8WsSEh5SgHG
NbBgko1Q7KaSE2/SDi2vWUNgLMH3cu2fsugDOJ1kL+Jao0ddj16s7U8olPzzOyUf
U1JaRC0OItj27clHyErQp90IaBuX2oDdM5vTmLXsMGaY2HG64XW/DAgMUrqlTE3U
C53MjIoSzRFJj6fOIiNT86tdJmLd19/N957qmLiZbLLyeJEJadE+wFYiMJrlnOcA
HObdyoijuecrFCilqBjNgi2dU3tfyUJNxQwKR4w5TYLlXEQ4YD+OZ9WMSF00g9Fd
r8ItRXfwuaG2Hl9FiAVVi7zK1YQ0rnPEQfscpoweaibn4LRD+SNDUKrtGHZqIHRC
EKSE3+cs8f8xgDLPILMZO9FnloaIfCHB02taOBJfDYf7VaUJ25FvcYef+FArPh5w
ZXu/Se2H+cX5rFVgPG20MpPRJV9P+cYny3hPx7citIUfD0uqVsMeibUQji/uIZI5
0PZKnYQAYW7xrrtPJzwbuzCmO+TEcxoxsmMtyPlSdX3F11PYshSxHy8xXrYgvV5G
uh4gWCv0X4ay8CKjXQFd1Y9TUUL/PtlC2Y2S0oA1EcNXM8ES+hJ5/rvCK8N5D7K8
KCrSk6rSoJI//VDcIpgfbuzX1na+Q/bHuu5W+ydopMORLrIE8TtS1RTDXsHa/cpV
UuSkyygtvjfQTlZXH2mhO7SmaSJi2TVajXTPsl5jl/LSswzYN7KQrEniZUbuSVkY
No4y6NbBat5Yda08Hw9c91J0meVJS8B2LQvTUPSBNOlfs2kUtOTRnOLRCx4H8u3R
giTI5DOKNoAjED0F1EkxgZYCnaf8MLD6AB35/qE1/0v6XGij0Lgd1uyWZdd2RnUF
6HJqKUdF0JPVIog1u2B/iASOn2gyeFVw33kibz7d/29KwU6uXAkLYj7usOuzMeHI
EO4KLG/3PYgyZfvOzVL9YQV1c6DrkBnhzIiIPk/TtOq0xJmpuupvLBXvvr2bVRwd
+KSTCttFllR7HHIKtinPQRHLNX0+gdospFwxf0emr0TmUCVfHO9W9DSPf5VDfDPG
Hd15l3aGU0NotwOSO11URCFG4n8Gtoy1MKSPMHNuupaXA1VxroqJmQrTdNu27auL
3gDYu07DptiKQpUkkgoC6kT2Fcurhbv408/Nv22wm9qI38tGG7HAgHPAEfZSxZ3i
f42PTqOb9ZUOqz9Thtj8esWweEJ+S1vrIAYmly7Pxp4lKkXjtjgTp02fzzeq31qq
XNtC/ojH/fZRWrQuWEsLMSlOXS55RvqIbAnUcA7DGb5iVg2gHQfU/AiduwM2UWYe
L9JYm+AOFZkAwZgAXE4RwA==
`pragma protect end_protected
