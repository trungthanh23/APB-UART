`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dpejivVhH87G+n2ctRjjrPG7Pzi1RODz69ce0/BQRsfs9IAjzoxrP7BxiJt+wI/Z
BSezXtWoAldF8qqJZDtZ81z0mrcCL9tgi2wSsckh17pqmt6EvYcW4Tm/KbJwZxrf
PaMJ9hBHlzBc+dr48+ChvPp4YOnR1jNDSNoJN+SZ3A4XchHTAuYMJv/HAN15MQK4
k7VvzswSeeQbPLo7P6eMxdDtXylajnzmNHIGwAuyah0vOG2T1jjFweDSqVfP1lxp
XyJ+97VzscZA2AsnHcR6XkQcNWdeHg4ADHp9+fFQtAm2UNMUSOKwsiTZ2Ku5tvhh
zB4Hr4GEJOd645o4GO6uFA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5312 )
`pragma protect data_block
zNRnKGe4IYTF/7ANuOoRLdG+z4SuvRbuHLRjKdlWfmYcdHQ/Cx4J01PgMCEyhebW
+k93OfY31nVrYi6zGktIeLXYF+uBv0q1irQhJSw2u+mXAFUg+NxfCxyPFLTVKncc
wOL2Ai3Ko6XWqJffaWRTFW8v8AXMr/iVIx2rb6mO4NZcJE6FXVI7U2ctntJOcSTh
I6SvQ79DyRh3H6xN5u7PMxRgvT47XvMKyB+slXaui0gqBvAm2WcQL68QX46eX1mE
75JYzBTOYltF936A7DS0/ZATqU/HJz0vGVwvspg+lSEbLANrcrU+rrxDsLQfInN0
mlueBUQwJ7EFVcoZUHkgPF0waJ/8foJzwP7bFWDzfyEXCq1M9DeCq3YNpYPtZ5s5
ne3M0xyvv21+LxsXScRd6uF9rjXX7Q+j9YTbqLvMBb2muj7Iae3agVG1fVuZmQ2s
353q2SIwcbxkakFZgTQ893qAg8h9qraaosEx0GlJiJahsi/bbYGWXDrZm5/oPAlE
QJML/Bk9sOTE3EgbL1ODUzg2qqT87l6dui1P3SFKOPLUwlXiPtKHCAzZxIqT+eSW
VBPhdtuyGnMYjYsylJTFMhb5B/pCExW0hWycWQe7PgDoziHpYggDV+a4uq7QXkLJ
uPi0nBs6esxjXc9VKi1nG33uIPxYj8CFEMrZYkdux4acWa2xxr0cBccklVRn4+x2
evoa5jD0QHO1xnlnII9k6WNya6RpBG7g9DGus2QKMDQET1u0zPvM6AvMKpMkm2m8
xY4qUlIiGeRbNxWNEMKs16sciF5IMQ3fib7fwEJXWEeqlKBEcz//eKYk+m12xhkn
/0gjFX0EFAh7Lv7njzF6+YeekzyPnxGfjHhyWY4vxN9STFow68kiLQW3up/x6qSm
jnuaJRPjEMO6qLbZPOEFdTN4vGSTT5vAxrZw3PC8nmnFUkK3+SvMZRyQrnTscG/c
qbRRE3QOETdqI/PJMEFYuvBNp6xfMVwQjrtyjyHGa3/zQBTjvd5D00ghcOzMtXwu
b0J2iSvjXgf4QQLZYxWeUYYVZpiubCfowccNcv0eLFttmAGpnOrN1kzfjKmnW1Dn
oCquLe0DFxR0sTQYotd/o0xtBsZsEIU2DziCLpGwwAHpy8ZtHjosGXiYvpj0YuOW
SYkYpRgxQSfuW121hWUYe/p8LFUaMlndTC/5DGVlaWGU161UnG12/XCzjiUIsnbC
xe9IVhs1rCYjT4N/CLA7lvxNw3HMYPoFOjs2pimxntAypNnDhJZ76wH/tt+yfgIx
zZLPZcDO+uTVwyS4A9lU9y4dbbD0bxVhe9xK2b4CghRYZkKp6YvVLst5E2qrC6yv
0xrzXO1ks6RnYvwrW6x+0cxvo0DaWTqcdQVBt8jZGYQyRWNWLXrfAoMfToWexfkx
7tNmJkqUPfZUirXny8ub+t1izRjw4fDMrS5X5gd6ydy62JdHq57FquX97SygTauJ
PAglsWCEvJH8oXKM13UVzJ7sY+Mpje8/faE5H21fDac4ylQmM2qS2EDevQa4pqTO
KubFoE1wfibzRN6Wnl/DTPFTOy65/WWMZZH2NxGuruqEZXqYJkd3H4xz7GWgudi+
lNVvif28Z5ipMl//K5F9j6WF6doThqgg1UnNumjAn9UeVNljGZHfswsFu7v0ftBC
5vQ7A7IfC3o9ZelCya9b+1zvk9xGeXa+GKk15WC8ZU2wYwVzit6tM4147Z4uJksk
pSgdYs/yZoEuId7NlCrueh7QxGIMXgdqyIQQkQmOFp3YAYeRlfACC8eT8zRVUCYe
XjJFnl5iyTUXPZ5oXyCIDDsN5GB06yf6unQAQc9sHJhZftKGBSX4dAPed7qP+Fh7
Tk3VvsqjDV3CzNAu6xX73ya0JQ5OYBVNq+Q1mWzhqo4OkDEejADHsdVuTMIOhAhw
TpQ+Djh/4A2+FEp0jlE+/POT8sc3P1u/RcWqOjXJPruq7aSKgyS/Umm+LX+WDEXd
dqnFBOguOQE9X5VoxUi9jL58qwcW1vAQAxP/TfrDNeLebWw81fVOHKVfHYCBM6iD
Mx26xTs5KRCMSYl9Yhm4pmO7AOVVXTtIAmYLpPKJ1c/M0bY4oGdELS7lmtkj4AvZ
en/WvFwiG20no+NjOoH3lV2puSaHddoHTxrq8LgQ8hpP2+RAS6KLM62aAJSTUHY5
FkMHGFu9iWsDM0KBTz72CvQFaX4daFhmh1/TNKNzOM4DeC6XUHrr4McNrREp3wIS
jM4jVhBubzr9zM0sg+FCvyHcTEEYZP33KUJD76fgO5kMZoYe3H1B69i7aBEUptfL
bdJkl2EW1NgkVoS/veq2yfoHrWMEk/MHNY9IMCNL8wCqmjFb7UOCsrJaN4+hLIL9
pZydEv9KUIV9djZIciOJ2q/jGCJYMHdJ79AKyjdI0dP0BBm7sNnE+Zv4P3GzpbfG
XmJup14DsrreTXMktpZb/t9kKvHmvegEejl6RNms5CaCkU5zhhyKWJmOhK3STFfO
rSAl8vrXQg3ySQ9+4QwRiTwzaDHjkeC/SfrZEfEkGVgNM69V1deFanoJzq1W7ndJ
7tAucBbkHnZLhQGH+0y7K7nv5h5birinbuv+vjKWT6lPthPN1SXUZ8f0GEV5dZ4V
A/ghH7ZSw6aZ9fBH+pv5RhtVps7nV9lRNpaOzUpmgzsKazEv3O7nnwczuLDZlaVb
CCqGQ7BpE17xsplCM9E1l0wdeh98fVSwlNNejy5rhAVywx/aa8THT5mFvMWH3QgR
/1AwQA6gOqXKmbOXimsAClQueH84r1m6rYRwUKRujr+E9K8Adb0ZY4hwSFZEXvYF
gDiuD5qAQfHlRTmWRAlsU8zIaiBd15ywsvZgIl/AmR5cUaLCia/UBFiSs/flgwCp
olCPDqWc5tpWwwCn4ASYuezFCb5wLrZBcKP4zCJpdws9cMRXtFtExPnQnvCanzBt
+1YW3ridV5e9mYmojsI5dU72/zn6dGVSed722XvbL2WHxS2HFKlY/2S2WI/pWLJ5
9GYNRYLZ9UtzjiepBGvKyHKIRNI/nlKxZG89DJc1+2llnb/uscl7EzrAZFHTPO+M
n+qOFc5mFNYSpaL8nv+qO9sAXuwNk3bJbORm63qKvjL2n+8G8fBLc8pKLGdB9Lk6
ge4oqpq1iQJnF/zWdjU9l3Rk4aY96Yc9gunqksZ9atbclq6dp6rdHTc7wnfbsE5A
5n9/3A+H8a9PJNLa/hUL2pQZ/B1aO80mGIRag/LuC1d3UhvrN8UP7HFBHvkRXuDa
yEgsjNv/RV+KzQ7xE1Sc/qwDWmUOUlEJjoCjNxZIc0g6m5ruSq/ca+FuHwfid+KD
nhO+Rc2agoWEX+BgukKvNwyNVppzEhrTEXwa+RSCaGvxShpuboeYqqxHuWWBZf++
RR7hvVmnwDYzEHfhd0G+nxmhaQZ4rnfEhfTS0vZcgeBZteqbSOJEGkvMrIXKKK18
D83M57LnQcsWWmq3PWtkMalAWE/mtN6Air4p8gjzIwcLsYjosmG9CfbU1hFDknZe
GVR4e22ZSxH1Zhqb4b4XFHF5kJq5lnw876+oCxewX+cEXW2dqXJzojerxC9TQ8tJ
yAYlBqO0rnWofFLzJPm3RILCOIr9gaDfl78lQBPyhi9AiWPgH5zFPSLxojO2GKkP
YtOC0VgEHmTsWgZWq734H+pwUlwOqMZZNyztETSURml2KOgpXmL3rwJkJZSJV+xg
7UxTzwnHkUS8ZlAOBXWyEfMVPigCXchGNe/8sNK2fsztswjG48sdpb8XjRIWFQ3J
AI+2PF7PdCosNrfC8Lztq2JFc6iNrA4qXB7jXw88iG1aTHHICShYdOeDBTi/FJ61
NeqkILhLM6dlpfOEwafaV/VtmSqqs1nboATPWS5tv3ueqHHkAFR71iwQ25KbWfkt
ZHVIE9FVGYzd5Vltl0rYr5emu3Rt5yToIj9E+tBtgnRJfYlJyvSY6NxtP04/QgQd
43864Tsci8+vXTtcFpgbgDmafM5iw9abxsM/NLvW3Tcx1a/hmpSEOVXlEl7GAXmz
bPjTHim6NMCAa5XnPNLOk4U7JLAp5jnVVwqXQMyj1SzpPW7oMAdalOF8Z9E+qTq9
uGYIt3yDnzjdisG1hRrRRhsY0Y1pZKmCWuAfeDxcdR8LF9YxrdryJvpdMGWTtskr
7ES4hsbhe0pd/gqhXxSov1NljVrg4UOIh0UTZ5R9fpTKFlJjyNOlRXghPRmoNbwY
c471tm8nUKm4iXsVexlKlpd/SlGzsrV1Q21MPa2OBvq177VErPgage5PumbC0jV3
TgpS6dRxx5fcGwDsqyHRqUKHxRRZIi0eKzycBL7denvYluOcXPdktg74IZoB0uWV
8vlj4m+HCiFBx7cG4TOO4uO8tMytraIk8C7vgMV49plfFxxdbnXVuIeBEvN/DbZm
ouMTS6yfk0ifV2ooK0K5y++As2GbotoEdK+//Zex71NHrUpV5uZJfz4kXXegn5Rx
J34xWj45YOO5YsnpwkhhM8oQ2re3hfjT/oLNALGKwfsqKbXYbcYMsg8/gKR9WAhR
FltiAd3QL6hySuHkk2dzOAxetQ+8c60Zs2+FKJE4TWt1H/ZFmXy5lSiPWxlEFoci
stgmBl41ynmOSaw81Td2CXNdED07cmNznSkFO+BIq3e2GutfT3wEFyDQPVPa4VF/
u1lKugwwCuDIWfSoeYiGbsNWF8tel4e+aCnCiz+Qw/P1/gUh5hzXw0FSwuqEUpTf
45SlC6svKszTeQTkSZPAtns42kvodjDlenxKLXw6BJ2dlDHJhb0vUhGSwDesNaiG
Vh/l9IlWHH3iymem7ES566rLfXMlMKaeo+2roBLTFbT9qGJNwNXPnO28ivcNyeIj
DQ+rknJZ7L/mJjA/LCjTKi5d1dyr2K9yIH/dhhLW+rWDkSwQj4ZiknOCTBnM955r
GFYZB0oxEBsf447xty82i81z0crKiFpXtu02UT98Ew8iGvIpXwjxVBbNoOdgYV8W
Ey8vrewV94x+uYQGRP0NPXpgbNY+VAAru9pCo+QWUisXDFFX+fXWLATlBaDDMK1M
wI1UzAm2XwLlUjhAonWaE5VwT4Y0woECmfrsRjnQqRZlx2x6BrfNdX/yaj0/zv4z
n17LKBctYIbumqWW3pAuETFPgNOGb9UcncQ/ik/6b5LOlA5GKg6bXML+sX7Vy+wu
XNaiwH+FJ9GqlogfEenSitFzUmgJEXZ8vAcDYbY0xCeychKlTI72CcNd2RB/Ex44
N2UiIoBb/18eWhtQRX0iCrnHj6lQRvk1KBCpP+bdfcxOJX7gdqaPA9Rvt8R5NsjC
waAJyGQ2/VGi27f/6eUElGK325UwsH6mhnrpFNPJ8MMB3I6o2KF7wBrSq/IrYEz5
g5tUFcPZj99MN2YZtAzodPfMBg6mp5EDeBPfi7ZMYSUwvDw6zMc3Bv3BOwbFt1bo
PuOrwRXj7k+wvC1cMziqCaM9j9wSgJcip9xbE4HN5TXYYpQnIrRJgTvs35ypWpx5
nxEl02w3vQl8k6sk0Jal3NH1lZ69sziUS40G7KsY60VOWy+rY48y8trU3jT/YIC/
fwmNpdg5qZAsTksSBSZ1z2UfXsa9lFFKkdYriIYT9F0d5A4tJGJBMXNhUEFFVHkR
FdV6ivw2OWuHJfJETUwfICjSaEYRLza6fVcAPofx4WPfaPFeB/z4TJHyfOfjyPI2
h/MA3Sm7AZ/ED2xh3fVLK4FaNy8rCz83kccDbxICdVDmAKxAykzkACBdme0FhdE6
jj2ragSBOmYa3HqIh9EZHBS8vU0OvJTsWz8Fy27jwsxN95Sc7/6LoENnRKq14LIa
lRSdqWGq5DjjSNBL5zKaPFZvoYxl1Th6CnGBP8sHaBTehkg+gDSkg2ec7/CxZZcQ
hNirYU0yWgucsRSz7hOjqwnxbCDbFPDVWdv9Sf0XhuDEKdfE6Le49wED6qUp3vul
XqEDjfiqO3882lkMgsKzK5ii34Cw/tSswjYScpoOp/AMO2h0nwlC0mwS/55ug+T+
BOGMMJjhXSg33ToBzsJ3qt4VF5t54mo+8ydnVOpQ2svzZ2YVsFZc/tl42HXrSwfQ
l74WJXB1iEs3TkRzlBiMuDn2u7x2jzTwEmy2ShYmlts+M0VDWuJ3wuDaRKEYrhQT
0J3S4+YTjDZTBc7KtOnklzuX9rTBE1FmzoOueKaIa88kwGjvSYsE9rZ2M1oynfjL
jw3qMpYBNcPczyuOFqeUpNwK38kzWNNZpB1e3XXposb+byi7rvJuGy5kpEU2+WqP
uF64y9x6g4bPbhQP80K4ylzmzdOPjiX51BNWsgZscUWPajdDl9FX5y1Ore37mwYB
/0U+iHsSUz7D76r/AO/rJwzQGkpsSneAo4OYAGyoaW/tQDyuMc/hXIBP5FhNMpnB
W+LTtIjDEnTR5Cf/CBBvZrC25EdxuusNFEd95NdAnN37ZEPlI6Y2yuRpDi3l5+Wx
8n+3TJTloDsmAO9VSFRKLWj9pQyPwZ9GNNdFTMhcgR32p+b0sY49Fop6xdcJi1wK
EsrqPAUtzfTS6jkahPb5iJ9nlKK3omTPNgF0Aoq8vglTVSXU02/2jeihfIXsQwvy
/M3OdMP8g5ZHztA9gOIcdK2YR5t9BypcQldVacI9JIOJ9d57VFqdmQxZThJuGh6t
Lku5yrhFE8PEwfmjIj+SpbLeh79LZ+AzsFt63icP4HgRzS3lzVfE6HF0lW9e5E0L
heGBOTbJSeO5D9jRMjzrRcgs8kty+I3FCbWar4nctEvSE3tjAbHYJYkLVlcvm0ki
Qc9ViSJ200c/P4vddgnYkVSDk6m3ITa8wqPzRHTFEjdU1IrD8sbZdYJ+22t6Iv3P
uuOytta7XUlj4u0R0PJDMBmOdwIiDZsKyZqWvMgfEnDv2506jFHIwHzvab/A57p9
jCixWku7VwU+YgxjmusXOtGHwgbfEjPHP1uo1jStDOAtRYc8bIJMFETo//5HA+21
lldM08xI2sB36kktCnJnfVc1H8sowN3CdGnFEtS92DC4wpp+YIBr+/D6ndR02RzY
0n/0TEwBqilR37muDWeyOqTYmlM0h4Xk03I0jX95fDo=
`pragma protect end_protected
