`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Zhu+ECJUQC2xncuGISoOJgpBXTJ8QIUipBLP/j9alsiTaT0EMiTl9GnvQe1On7YV
qJKWywXgCzvCTsMKXUGlTtOtk9jn5DksSUAwQ8vAOHejlEApcHbLIQts9HZBLO0o
plCgdZU5dLL5g912QUgsGqhK9nJiH+w/HJeCCmhnwo94OFzo9QW7mIFsXf0ufD5w
MLoQ1G+xHy5pyA1s4cIxENzTs0WDkckFCjHMnkdPV2XLpkBETITiSQr2LiTDZ1ZS
z4iB1WtNQsrXZi+3sXY0qpTCnlap7lv69Hv+5qsDMuGhYIlh92FtxrsahzN83KR7
2OEhqrnx0YKjgUlE3GRzfA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1744 )
`pragma protect data_block
ls7zIVIQ7n6x0AOOskM0QlmAm5Dam9Ib2zxrFQegN4ZkUYGt+WhNIIR2xh3zjtft
xvXejoVl4R2XozSeWDntFkYSfK1e9p1JlXbgHI/ieYVtCyQp7RXjSxP4oHiQ5V3k
rRvwYY4WJftFB+VSmFosRJghB5h3V1Fo5EPoUmaAgHSCmcHK8exiiYoFsiVWuWrD
qDXPrs0wKp4QnsUbMCjTsCHSjUDAFgcQ8UNQf7CAAWVCPyi6T3kv0IlGPvjShIic
FfJQwoJXI6/8FCbpFA/86f8st7x2soxI3r3PutgpPnSUo6EzETbyXPPkvPWUAEgu
UtYbVBOdA02x3w0wQhwbKBoJqs4zeaUkzK74IlocrQ+Si9AlLILSYmNtEgXV7uj5
50r12441XcnXz0mq8fCjOM16mEtFjuusDCtHMQ0vOYTR4IUZLWUdUsDCpBEbCBs4
R7konMnSyN4jT6N7rt9N0DdE8956UGkpTB7gii8URjlcX/l4M9zNm99ggWd7fLVK
vVVMBDaIHk36IRKa/wFRM63ZBXYyUCKZrHcxs7LuM+MHHDby5tH2GXvv9egAQg3Q
vhlahVhgnvnS1pcxZzJCQRFyOk5ALn+pcsgYjVVFBalx6Z1BXb5+AvjD+rMGDNnj
T0ZWV3ANemTBdCfzy14yDRWnwQ2LRPTYhhHapGMjg2XsY9n7VN5ieYeNB2yYO3FV
FCA2aSD0o5SGbRsHJ7+kBECSdn7/aWnSTg9xZQdcrzwI0CAcD4EjI5Wmu5KHr3L1
DGzSrjEz63LMqqqxOqFMoPHR3Xe09zwRzldoPzcDt6WHqK9fS+KDVxP6DjzO/wE3
+o8HaM/Vd1JZCOB7+ZB7xiaZcvM7gfBZl/4lFh0D7xwU56TQ/TEp5dU07AxMtePC
hPOvSSmnjWSdobYpnF3xp4WWwZy3oqpYLjIGEiPRM4tDB9RPoQIiUD8+5dzstn+e
XJp+/w1jmGFdcNgy4y4/FOoGccpHUoPq5gmqM96FgfBOv0M4+jOc+bwQCaUXMPcz
lX9Bo00Fy8JvV2RvfwuS6AsBYUNO2+t9MO1d8Yt/3AHz8+AGaIy3KiTFOTKTmZH6
3b9BpOLZSiFBJL1I4X0Mx1W5CGrnqd5EKGNa1bjU4V+QKhsHTMy4EBVrnXPSYa0G
Lw8gjXlPoAeykZ31pXOWidEIs87HgA4/dBfp1wrtGtDCSk/J/o7qzDWJYUek9ff9
9bSx8PWPcdsTvABi5u2tPHupGECSb18P1voUQXureTCWsnAISRbRBNWqJdTMoOxl
cKK9sUQkQlYNgabQoVs3Bl784JaM/eQmhhAjf1VQq3GWOh3nt2IvheLOpIvUx6H+
2KuyQcqBHWdlwGW4+q9YhSkGGDYmYyMeWSTT4WrmC6/asH8m5eXmcG5kuLnSvXgH
1rqrZa6fRb/qUIpOm1//+Wf0yeGXUmW4YIwQviaOrF9e5/hEDA1WssY1b5haHz1V
kx/CUlOzpf7ZYDYlQ56I5oc832KCkAO94UW26Q6t/HSt7FvLToQedNx9737jsDnV
RaRhNIB56bR4IVTJofo/sD/5TrkeQiIf1KE3fCfNzl8GWXQCLSgbN94lQ04nnlv8
qpS6/NbZ3r/GIobWE9g8IlTpbGqTVgftt1bTr3dwfU9qUUnLQLYoCc8KId4Oq0lm
0I9MbDRqbRytJDIdewx4oC09+PlmEZLSY4wyyl15JJlteIlzkeYMgNRHkuMKYakG
JhyDRx1v6RhujG8p4GoEg5GTB1OFBYTNfLhDDnP2ofo6LDRo+sUPkHZa+WVENPph
kF8FXfW2BGhyPoXPWPChQ5Yph8JWIxGPIiI4+JoLz4V5IQ9ozih+tibE7t72yumR
qnHgYYjM6WijBAqnKcUaPl2NJqnrO2OpKWz1hDnzUE/Z3JVVNTJb+X1dj9gcGpkZ
0FBTeg0niH6c55SqK2ql73tLPmt9uGjlLkASF4cIg5GKVzYKu8+jQK9c7eOOtUDw
eM9m2JUr5961yYnY1Bi7ME14t0V/qBC6FlUvn0tVtf0bGBxE3DK4MudV5Xa0riKp
EIlqUtsJlRVipcLtiGLoA8vws8dw2XQrqIlJPzzwUIyXEl/TahSyIDMxvHx/B59+
nciPmnuEkjoVlseAf5v/fDE1ghhGVoa7hJ9ZKJz4jT2utmxeqNVAycUel0+dBVOc
vOdiL/VI9K/39n8BkCyVkFfqWhCjldtW4gySCcO8c3cVFT8v+W2bSN2cqlDZo9Xm
Kk9fCm4GxlDrQ1Wo+iWaqG+nubsmSHY2jJ5xyOmyGRw1yu/lCR7OmId1v56cZUDz
CkMLuPxBNh+c7sOsc8lRcQ==
`pragma protect end_protected
