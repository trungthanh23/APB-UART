`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
h9hMwXHjbhg5s0WimCbR+vOW5F6ajCsY2WbljOPT0A/20HcuUPWAZhqLBMhN9u3U
r+B9aKrSoh6AvKzySG2mJ06YG4Po9a66GOD9tQ7KNcfXSFdSUNCTrnPM6M7eGl/S
o7FSUEewuhceQfekxbnkpJQnhr+tXPGkxr6F9TuMqx+h7rWYN9REKGgtvwnyulEN
y8a7UUry3QevnSvwwrEutU73xHGbK7L12kAni3+nYLLvbjLEWuaOKnG8hw1lq5uY
uvYve8t8mDNIwVKXLhixyLj8mGOp1HJtu4aWb685F2xZnzE6LrnbApDANFIhfW0K
e7vXE1mb1U41jNVZgnsNYw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1616 )
`pragma protect data_block
mg8ax1AMBSBvXT0vHOiITPpdHNmZGPGWblZSC/OZR2pEZhYpoS5gzdjZrwZ609q1
oxh0eS0SfMb7Kw93nOOr4LoVS1JjcaHFMwvgNPPIJzwCdnzvuWdAZGlPj2AHheDt
bX/KMWad63Hj5Qxu9t/lTar068H24EUy8mqfEDbPdiEXKPr0zqNurgbDCFcnQXR9
CUDZTF1tntfqF/dNv1bLCPOWBr1W4/7agsEUzMv0E17FTHt2Sh0g09HVvDJNBjeE
PuAAUbERAZBU51+17Y8WI7w+FKbZucldKr6k4us1UMBNGuqNGmEvBDJ7VGQ3mOuS
sZKlfH57jIzQ4bD8ops+qzwJU3uzX4bbjBT6FWC2KrBXG2igQi/V05XxE22rLwqE
7YFlsgRT8cQnWekUmEoh2saiZ+FAI04P0B2DExDKOyZCM//WYexYM9Pr/2XtbECa
h2zctcXIZztcUryLQ1SX73Z97C2olM950KKdbJl6EGF0wkVYcpdObEzINXAgqc6X
25B0pIT/xHMs5ZUJC1rTGcWWJYT8MQyetGbIAK3UJnhavOqEj6qtgavLy7aR4hhU
Z2UfFbFQbk7WbOeRdP4WNT1IlXTWEW+xvEW6zHzboRpDRIC67vyWMICBaKFF5L5v
E5jHZ7o+N1PWHkpN+vee2DrB0HdAs9WbI6i5fYvIDQZEHRxQONqj0FWQ2r2Ule4w
+OxVqZGMgMP8rlkTdNno/IW2J61xMcR0XzM3+REvGzWHmuBs3F+dOVkXLnfH4B4d
YysnFOPjqhh12NkfyrX8To+j9jrrCLJ0hN/VyKv2oUgkIReZCYVUUzRBxPyOCYPn
9P1VriFAc7prOYR7CPjUGR0NoffpT2pvIHJcyaef5lYGgePZ4rGrd7mCt4Zn99Zt
V+1F32eroq7lxGaVvt0An+nCc0KnjF972sIwikXRv6pVQ0PHOLQ9fBUmS46nVd4m
62wZeRGxstrcUjg1/5+YYwMC2U1fxfzaofur6rYcLwptTTrIU9Sq1jwbjjmfsbeX
QxENUH60m8dUBtkv0hxYoDZ3yz7gDPr0EBQ7O4fGq9KjC/1RmrEoJT9YH2Sgxts3
wnOKoONPFSu4XwoaR6mgXFCdyRVPx9XYEGz7Mw4cFSfBIO/BgyuKMr5iS3Zsn3Ih
t5BMGNZFkJmLVThHabD4nTAcmtiEfiKPBOJeGNi8kvupeIUZteKbHrkADJoPuCfX
cTLmL5WGuDrWE2oOQl9pwoIj1WZhkOhm3Wp/z6TK1FLe35WgC9/m0V8yH3tng7Cw
KZzI/ADR+yULK1M6UvtbcOn+6TASRLgvDX8v6uhBZIMreksJryc+Fl47hHQzJWxk
u/fuGl3e3A0PbwABSF17BrP0nuI14Oug/HI2XtQtQ0Eq2qhE663TpF4TmZfPGzY5
VGPnjIEko+RqogFjTCIK2aRkHB2AAx5V/t7nanCRwRInL30T/gyt5rvR9XrYYqZV
z4G/FCvsdGca6P3sZ+yTyEjqpT7N44F+DSYDDQnkoSU9py+AURW3/mVEAzdXxWSR
PnjEVTP9LIPc3m/A3yxKxWepHjCTgp+jFnlxI0IqHoyjvfg/G4l0enZEvGgX8cTE
IKXr60IROdOtuXX4/4M4wnvOaN01e7mhQ2pnAIfmO7BfpcKSxWU/m3WegLnyDyPw
j1DxTZgauKGS7oSgiuTFISbEqbReVqax8hsC+f9u8yS/gE9rqvabeDyI9bNuo6Rm
n2O048/ivfJ65edl20evrKVhzF4uHpLf0jSuqKrjdGM3X8ojeQ/ZwE6bmpqWL2Ka
sesiWTYUw2zBqouUw9LRaWSz8spngFo/Mdblg0claWB3VsxkHNGuffrNmYSA4zpz
RgTiuImPbNHAfxHwoNvUdLrgZT7vwnvRgn0fzJypf6BiWtplYomz8XHSR9Vv0ujE
IuMB9A4ApH4jbfHVmlWYw/s0+1EGb/EVsk6DkEBL4ZBeQlgnw9esLqtBbfmNlqCD
B0emoUWAsVJ940bruf3hMwr9IfpW5eejP2J66wv8xbVH7ZXL5vh3f6mzlKGP60g/
oxnMXlAsVfABrXJms8tj+l6MCsd0CCzt2AgQO7IxRX+MgCkL3p4okW1q3wmmB4tG
hrqiz0uusUy1mMxy+C+2SqD01AKtgg52/Fq5pL7ebcc=
`pragma protect end_protected
