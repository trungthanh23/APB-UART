`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HvOFIdb6gO34xEVPwHRSDkSIRxGleMaxgxy+xcuzSVqMIvUTu++ogRAMb7D95NFD
FR+YcYqKyx9OdHLacqIyXTiS+r54jpnzbEoZV0G5JhYQEdrwufL3KvJCw926++9A
XfQ1GlhFixAwsP/6r+WVRwUz2CS4BLvyT5/76mjNvyhOcBDcJuytc37D46C5i84n
ptsktBukRZ9POtvP0pvfMURg56zHaf6C2vpsC9VJvAlgEReW6K8VRRkulcXwgZ5y
YgoGtyVYWFpiyg7YLA9xhugGP942QtbHd5GuAQBu3kLmxBzb2aTSqoFSdyxX9m3p
As4RWKXp7osf0eKyWNtWVw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2224 )
`pragma protect data_block
ktvugRoG2nDyeixSJlSeqZgiYjIaXrMW+g6aLDH1iTf2YzDMyEsGIjiGNfwC/1Ul
nW4VGyzzb0OAs2IeOBY0RO/4FKzzU0be7lTaTdelBZUnCBPkBsFz9pBfuCalxtZn
H2/71fcJVTDPD0haLPrdk/sxClsTW+aLamOVAotawGCGTQ8RS8Nxk0RYwhzO8xZK
qHj35HXKexJebIQwsHhnJR5cs2uPru7+q2inIcVULpE0dXjYhfDSCwBzS8fpPM54
xm7VaAefZ0Y1a/Z9XYYkXWF6V5qTeo9KFGMkhbLNt7Tl1RhvbFXOlVxgyOkgazXP
HS9hWRWj7ykmMVLGeNNJJSiACjpA3iyW3Zullu89n666erY4/TX9+Kt3H8BaQVqW
QGk1B4Gp3pLXFpF6VcTahJjisDuuRetz2SpC+gMeRgs/VxX0p7m4hSSjLCjdbQlJ
M5WkCwxJg48SbFvkPhpOpx3xD4SSH+jDwyrM/zsbVfEUJOQfN5TxFpnbPGDqDhHo
X3z/QJeYI1rnFfSAx0WlDfTp2Mo3Aa83ulmdXK2fh2czgKbgRefisUbSUYfwYKGQ
EpDwhg5txspocve6uc6Jri7uXFiuzJfg9DoRpx80MO/J3PGhxbjitz5F6pvO+YC7
tOqSX16ZFuf+2bjvMfVzz3Ihwy5ZfgtKHGe7bq+1tWRnsa/K6/Ew88+kj35wlTLM
H1yjrS/xq9UGKo/PpBknmwUeuLc3EO8b5uLHszxTViCBEMztdwUzlBddPtDT6Krt
hrsPJNTpMb3glgzued9CXFGjm2k//AHmjXgmYH/WZ19Xy6aaB6ZC5pr7C/S2UOr7
GBICkBFkg/d04X6t3OnaP7XomkztDXMFecLdLUIPRpmgzgG7ZsqxsSj/rToayHRd
eDuzysYaU1mZfezW0BVZrqTrTHL4mkUfE6gGq7FmxvlZkv2BNkzgpRg7C1HF3Tv3
jhr5fbVk9CJQT6IEDRU7t6NGY5lsbx/7JOSO4Ah/S1y1YCKXs1q1TKwH+bTFfiL4
4hgepRDzfBshaU3skvKA1ZVILnObhqpxFsk8qiN2djiX2K60TVobR+9USNlbPKeq
wo260jO5SFEhveSf+oGwuFS/QYY3tSZJVwuYj0+/q2u3FMKp1cGCQfMeSDkxBhYs
XbqQEhs5gYKCAd7xJxGwW4AUaOBEDohafqAnoQ05GhrliZ0UA6LwaaaFwiMzgj4F
Uk8jDFwFXedgv7IFjBr+GwW76ozVIcR9nH02xCRy3WxpfLpnLdafVBWido5F7eg4
OeHNf/ohvizjlJ8UJCX8yReU+Kx7zhKHK3qaFdI/v0Rxi2ckcQ5waVBO76ru5wsi
L+6jIK3L49XYO9vNh8kOyAT3B04FepVmN9+HKqWkjAJQvUs7gKcELxX+Cik3E3a4
1Qifcax5hSCN71LgPpR+OmGY5DJSr/cjEbRImrRQ0vScoAS/6iqwcAeEEe5qI4Mb
XipKynGmtNOlaGlNw9J/UedA49DQadEt1CUhJ8KXrp5NJNKrpdXucEI03cQMUsXx
h+Ps7Ebk7ujgOgBbQYyTXMG5Vzd0Exh4Vwzb5Y0OjxuNygGLj8Pmq7uYUnIww+nc
D8AQ6KwjdzYi/rP71vvACkALNOIujEOVHxwy9MZUux/xy6ulUmX8qKk6uigk0aGK
5I9AlNFKuKfYBK2xmrZK9r92Q2PsK1xsb5auq4p3CGRjNKvfppnWccGKJkTJtIdo
+deiCx07LAW64PtEZIInKOEhOXV2Ms1snq67oDd0neqx+Yw8pmsilJzsXQ4FLmjR
VWAue5DtmlgiqYub1GUxzyBg0ApGsMmL947udTZO/yX94bjBVeKCAB8XyXCy/7kW
wgSZ4zIUtx3nFWHbMRmbHZEh1TCxzTaWb7+D4iuqdzyjNY0zXUnDP382kANr+C4z
w8xikotHjAkjcp3GyBrCBBjgajEs9+/hbuJvjnSTE52TJwc9zpoW72puMiHVpHtk
nGyOyB6Y+Ix1D0efdoBQWxWWkjBPNYVOx2YhCHZl8/PVs6ipSYWX+2oOgey0N4t4
LWDyz46Y0UJhlcHOinDeB83xs+PO94Tj55+mUCUO3vb/ZHN9uqaWdBhQdX79YVtJ
fF9Erxmhuiuzg9+WKxs8nlACqAEdiqYaw0szVfn+j4UffLlph9QYrCRNDhQJ/Vo6
oLAjQTI/MvSKgp34mbY+ptmAWWuxs5hJahfd3Czgm3SSJ9SbUQyUAbItG14/YdpP
24AFdVLl5JT8QY2Mcl4gLlNPJNsszAnuB+7/ZfwiX7J7LNoP9fm5D+D/3YESxAOx
W8VuQrs31Ac3BSnBPqRRnpqi7NvfS0e0SqoauzmR6I5usoWG+vLNsWShGgmxozaz
PTl0UEv/Gm3gzhd91FmVPgO6F8T7qH25UhmNOjO91V2ciQvLh7Vj9pIx+gTKx02G
g36RpZmNBdMyDy4xAE8Ab7U3SpGwUUdbOualbP8IM3S2dOseOw37NftLpswOhZbs
swzDbBreAgen4qw2PhCCNrksj74hcecImQ+YGt8i4tsJNpDa4iHvbt0ClGjyLUnv
Q5sfWpJxNNkBUO+HaHwMu6azSjNq1xnk/lU/eAigg3xiYnS7YRKy9HkDJSZwFr84
V3+ylCUyfieefzQD62Ltnm9I4/XLu9/8eWXeH6HK3xlMhvksqmXohSrJfpuT/dj7
ErTJau6Hj2GeS2pKyIbp0aJmWNueJJWRNZdgiIJ31YsxiMu3TviQb9QQtlmE+XzW
NVmpEvXrF4Z6Da7A3+W1tUmETvkZdQ+QwQ7rtY2fX5ukpn8xvmvtMUxl/Q6c+fTH
4lgibw35Gl9KIg1p+LPfrGFqeM+CTnNwjzCOOfwjvGRdY06TeYOlV61LpcB1rBP6
WUrHcPgXuzU2dNyPYmKkOsoQ4zoHxi17BagHOpFj1vbeCcaxKmyqi9SwA1ZXuOPB
neoPJOAnI+IrrOYtbJNH1g==
`pragma protect end_protected
