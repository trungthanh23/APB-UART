`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EkzU3f2HdwtaK5bg/hjbfVVWyN+XYzTE4pGzeIC1hkpFWIXhyTn4FfSqhHU7e/Tz
jVLye5X7eI7kzVgBpAuGW39UnV3u41ZPqEmt0u40WL99W4krtw/DlSEAEMgUBUqT
bDIIWUmEMn0ArQ+RyK4kdNDvH+w3HKhd6mRiUG3aBFJZu6tesxtjT02KMi8u0ahs
65ySHC66GgDggLQehkS8CrHXqaRMgRB+Wx7CFRjcg/UJPBLG05+NEPuawI/IZUFb
9dT+WSV6xkFuF4fkPBXPr2zgIg8SsYm0rIEuYmTPT7ZUHFm3BegifIFPeQBtr+pW
BAOi6itol0LJCBnmGVDwnQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
xHSnw8qBSGe6LelN5fVRXhmFYnj+xx8sfb583hk392mbRgn7grYWLdj7Thl35kZ+
1FCPehEAWEqOsCNs7eHpAU0CxfLCoIgNU7vztD1UEsw4QwAIaI0iFrtsEGrI8YGV
PaKSL+p9SOSJ96GpAKyNAqTk5fqFqNv7QCsCxPnFgONAqE57Jb3S0BVVdxKvHUbl
7dHpgOW7BDDMscjfBcHyIZWH/YVqL3Mx2eOiTHwZsSsB4geU47B1NCCmeR6UdULV
cVGaMNfPTvCm5KS0cVOwpB0+I/GzPkjNp0HnL669p0ZhlGT7653vHQJuYui6ediK
P3mSXOgzsVPmeGsIvaTXhVky6UWa0RGOaAyR8tBeU9Cgx3cJHLQYTl2FetyN4NKh
wSOy5XofHCKW7gCucJM7TnlAQo1zHAWfRavI1/7CpWnPvtEUSbjc+ButGRR2d2m1
ov7vdvx9QF7ya4AntFzZLT68T1Bk1JfU/hTKOcsvktoWfQOLkvBCdUvuBuIVcsgC
AC1fJudtaZCdUya7YxZjRSkqTLUIEIGNJu4KKwAd6cSy7QSKifU3bbQmSqltVTKy
CQ9TtH/OS67AW1me8hytq5jpsR0ZhwXhTmOWwaHRNcXksrLsWFhCjioxwPnGRAuw
bZEsnY5UBnBjV175QkIhqu/Cl32PSiTHWFZEtKxPcHRDseeskJJCfjGjijTbMarR
7Zw0tSK/oNAQMy9+u9tmvpFp2Sm1VSvCnl9Fo4GhoZuZ8pDBndlq6woWrt5DNlas
jM2rrDFkj/7OXcClp/TdVTtUeD5GDydOUay8WW3j+kqRu+pIyT2ktsGMK37qjEw1
kzGwUhPMNbINcBtWbYqThmQG9e7iiRg5r+7+wb66hzPrVDQQ/2oDZKL51sOE6WT+
+3U8N4lXU7ohOtUS5LLmvC2j1TO3JLf2Klu4Mz/9K4O5/psD/tamlkwWXj1GUMgC
ejPpb7LzcVO4W9IkrQxYPLWh0IWsJBcSFR91jo8YojaerJcFRUd4NhKYqXMKSzOd
xkR6D/SCo0f09UjWYUjSnAewGGnkqMch03S0VRj1d71fK2wMUMf3PgCtPRBvfE3n
MCFYDDDQ1XExcdYGuITqbvNMFvuyG6697lB8yRc+HicGX7Tzsx3BaVaDDgLFqsvt
bvEO5RiTWSJElY82HU7a/mHaTmXclQNJKAnZ6+8IOhdAril6xUBtEYhCCdBsuPV/
9kBzaNBSXnENAQPaxehTTqnwDUATyfZyBflLqGMfG2OKWPieBOoCpC4jOwODCT3a
lhmDxPw7xHZWI+PZ7g3PK+6xTxbLROftmzdCpamd5uRfu1g6iNuHafBQAUQRhXuW
eqCPNnlI3cXEdC4PPfZlSmmksiSmLzzcoOIeDoJawx1I4PXwfM9tbeipk9t28qWn
J6Yl9fi4Luor4mDRaC5KK9gqtKHmotBiohc1z70Th/yQ/59s66asl4ANNHzzKz4V
iDIDOAzn7dDsBBmcCduucsiU3sJZLzrjFFubVaeY/5GBxnwTjdwo5lS/sim2w3dS
Vl7KRmb3E+gBvK5ri+LkpEC/WJHPZ6dgpVoqKF9oq6ymhGyt4b+n9oiUNDjjtDEK
mldSwIyFHVw+PE9DpQPU3NdGakmdUsasCLmGynTxBkcafWejaZgv/PG6oTHM6Vog
N3wp0hHO8H5k0QU3up2cyMT8x0WhtTWpc/UtLTLPHCtDr0UuBlgVky54PXZ59Xa5
M7FFrdanksQ1JAkIJsCnHyNW+CPnvSYryXh+LOn/w0gXReeLnIMd1RfPGH67BV7+
M70EB/TMJwZN2WSj+0J3ISG80RpyPgX3zR+dL3xcHBPoXAI6oL6ZKO7KQ6lW2v62
sEFOqNfD5L8zhChRAzPmpip7P4PETZKYcAdFZb5uvA4E3JklnD6qSVBRE6OQPjw8
U5FavMW9v6V2IMuCsou7oCwWWEfN8Zu7nZKPxTJuyCw/HQFaSB98+DswCx4igzwf
SAkixifvf80nDQb21kqstqPimoCPsRCdxrIWWNh0qCs0sHYSoung24869t+guALb
dOgim+WRzlER9LyVB//tOCP/VTzmDZ0QTqwXZLmJ3NIVB9zudmAJY+gEfoDhRumn
XLUpTnWLSH6pcUk7SRZCm0DBkyKAa0npT2DoMwEQwFr+u+A11lNY6taGihLm/14T
38hCpBsNfCyrUolDFEvhooWkXhMPn/FZh884+qZu0SoGjM7IB0vHzAo9uUyAtYOR
V2IoyTXKuDYFiyEJIcAbeORK2cnO2rCpuv45XLO33qsWLpz9JrtMbm5cmzH7hDWm
jqCuiF3MaM04sPJ5muZlz1QDeiBbRdestaPx9yqXvrBkX2PE44tuvY7mfVNeOyRB
nO4hXwGZ7rf/QLsMusg/WQ==
`pragma protect end_protected
