`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
q0lsZ51oDLUHKqmReNH/1XiGQL1o7WfcwHiEU7HTTdQnPeLkXoaDYzsZjla3/H5s
TS0tL/509hVQUJGTWPoLc5tvgCYBx+1gvogBBVojz2Z7BbQ7W4V1wFGW/KVoloeI
Oznz+zfJxbIvB/hwVlTmDvmrKN9l+Z3SISA0H9lC3ePQCiegVKdN292bKNXk+Ck3
t2qJ/filzwQNx3cXe0I1kjT1I2LJyi3E2IPhy4IJSW32kOM6yAg4QMbNyGwaOLWJ
+kKtSI/YwpNhynbnpruF5zrcq7yRj6zrsSqTucBfDXCiX3qdyNe+ZeeypgP1vuwr
xmv/kS3emRoBOFBVZ3BT2Q==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 944 )
`pragma protect data_block
TGQAtxGRVY8yDXlcA2JAlAdjLWnjl1n+W+45D1St5+7Jq09z9gkCu/wJP7Hj8p4p
/bp+7133f32Ei5gbSnpvHge85nb2VfF9BuFS7WpqMJJEciYicRrIyUVkZ/mZGTTV
sISlUCF1zqDOcQU50c2NVW3hyGgsgxjIb+1oOhNVluhbO9Sq5CMBfCKxU7JDZRhI
GNOZyYHYim/q28sNCnCgZYZVwwsZIaEhF4OgcS4DBODWhuqUsRok1XOa9SnvpfJm
zsaTfbh659WJwWsdboH4h4K/J2ukuK3pqfqKZiTytyDdJ8K5QD9EWqu1tmHT9KJq
zmkXx12UB+d7LK82Od5ZGqIhXhuMuUq97LlTiSZBFv9rk4xHLjRA6Q4DmOBb9/f3
70G2MLXGzOeVLmiE9f0Pl5HMkO+/tc4UiLL8uBRo1IwINT6fhg+YI7K0bLV6N3QF
q1qhOAaJLL+DXEmLzltb98WBGvD9uTlCdju5KD6fZHv+5nUa8X6bMuxEybmEa4S1
Kji/riZbqANK0lE0c8XyR8hzhx1hrFzJxHyjBs0EU18XJpOHIjPN1cqkKaCe8by3
DElC16Z3tT0eyDJuc08ZWbw/tQvBsjGiS36+638j3Qp/d+I1Dfa3Mbo/7TPQdcI0
7oMCq8erq0TXm3DSIPuBRyj1pDyhVe4OyUiNSPGrl4WqX6JVT/csFngzJsNmeL/M
/uR4HR4tgNfqLx4xNEnJ9+BNrquP1Eh25F+l1Kl168KWT6y2r+zmNei1KJM0E8zL
8xk9rM5Zdafkyg2wUU+rXC6gDzYqPuk7ZF6LP8WYnvm+XYtfUnE+8S5ugJw094c/
8upGdF15OOG6x99CNwwPIboglnkrk3H7aWP1F8+1yz38FU2WC+yz+E7KsJjlPTxi
vpVGzZj90C/im9aim2jq4+P8/mJC5R3USRwRnsUJcu473rf5ZRXKMdnMo60GMtSa
KTOiX42iySyIFbpSfSG6QgcVJp6wQS8mHkeGrzxj/g9UjWgaOQ595jLTIqDIWdvz
RPXwNmPuft5vGOceg+REeSYtPun3bU/s/Zwlcxq3C7Y/r+6QlABMGiFRftnK2a0u
FS3psXNQRSCp92+EpGIF0bHqNBX1MjqqRs8VMjLQ8CKhs1igl5G4vW3vSuKziYiQ
8KLxRN/9p/MfYJsBBpf6rmsDSqm201bmwHIO2ll6Ea1TDR3iRMwVDXNhdlrcqmGi
5jctqYFcZDX76Ri6e5Iwbe3SRRaHQQYYUWZO/sNuTT0=
`pragma protect end_protected
