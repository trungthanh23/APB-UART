`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PynF7pDKr0f2RkZmM0ao5wizGSlpmCUxewg8FQEywn34/Fun9rdBrxw0POyTSZB/
1mv0d5S7txCwkMQSmBNjkbQRB5E0vYi3oCWSHT3HJFvXSbkG2ia1qhhxceS9V2B5
A/QyUTJPGchf0ubVYybTWcP6PLd4L6D9UxkxMdl68NQEAM9r2QqATKlXfL0HxKSt
3Qr/mIfXM/GcblxuUU3Cw/lUJpt8WiWQCj1kw2lgiE9YVwovvnOF3qiZ4SBn0/uB
gOzC8pJdPo70qHLqX7VSChoAVPLOUq2KgcqAybijFYX/ctuG01UFq6PebmlKFDFy
dyZYR+70G7STpd8PwSsCIw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2848 )
`pragma protect data_block
xuTPaiC6A8Ti3mqHVyMdUgRHlIWHNFkObcYrAGY2Tx34Mw0l22ywRIQMoiRSdzTU
5/3ygGiNYJ6BH/i2Pruw1GVIQwhJvEdtwl1yZ/Uab0RkdJS27d+M0eWhFIH4nktd
wJtWE5TChB5rMllEgVrOa/I6EFa7LHVsBvINTCPGKzwnTXYaLsl6ZewppaFKrn+2
FTnsdwCXdT12HWB6i0xUbOSLFxm0rr7PXLLy6r5R7pDeDOB3a4eFXmMtiWw+b5WQ
ivlFDVkyyxBVOFEAtLYEMGdIit0NmyGRCGm2bXOZooOgXnW+G5ttHOMA4gXp74RW
HUigusqoAc9586qQZ19ADISeCeb614PachIYNdTjIHhfDQiCHIMSXdC+cnm+lDaf
PTx1ZmERNpqYDDE3keSGCmX7L9eHK+1uf0OLR1lEVkB6Qppj0/hnEgWCNlnarbj0
79oNHMAu7KfC6XeRsL5urm0+jxQqbq7OIEohz+gWNn2bK4W7LCxeyXE61frIPLbW
oPUB/zA8CU/BQ0Mulf56jKxFFzw/43RwNtka4VvTb8NGlyNDhVLOjPHQpq/UbG//
TW5xDLqXDF4QKftnibQD21tK2VdNdP6yRTQd4uJHIZ4jgS794uVu1/VCVWylE+LI
+46uk55lY0zPa2hc8daYNg0h2SSTLHVu71hkMfKBujd5/697bVEHzz0tsEWQVHeE
u8lyg3k/HBXVAAkNHH09Q5VUeooOVmCns8ourLpe58d26qo9krPQ9tei69eX3dZ0
3vxxHyJxLyas9NyDW/V7kbsEyHe6e3PbU7Z+bFOuc9nXinqYrCpACaxihSWkw66l
DpafAENQJxJapoGd+lkf0FOAvXOj0GzUKMCa8UnvZONOAN4ZLoRHZtV/tprF/l/k
7/h5XNukUBVrRSHNeNim7wpxvKwA8j7QKOF/pibrgDczOoF9VaJDILcF3wZwQwgc
wO5tIfVd7dbP1xYPXje8cNm7f49sTH0hSg04jw3Meix/NQ7PufgWMh5ATFsbnefk
nHQbRhxbmF2V3PK0xKavaUBMjmNEuQeCtRUADAeFD/0+x15vbC0y4E1VTHdPVuTj
QdLTDLm+DEShfghTheumRiE1+/owMPyhd78pOqCJzGq9KR/d56rXjkhsfynt2cPF
hzF334R2tE3FOlIF2Q/R5SjD12JSBZPw9TW/Vs9NpHqhhzBbcIxIXLXmEPtlB10I
tw/L+A5fIOhSMtbHLIOu+zCHN/lnwVkSohF5Ru6Q2Q1vcb7zpjZaVfgnqGmxwPk9
UVzFx6cmeg7iDiayDHQPfhVlSNKBxcrVQYPb96ZKzNpRi5sRD3JUH73nXDZ2FXVI
dZQHvhvi2oLmzepY1JGUo3WlVcb8911EO/qr5Uts6CNMrYF8x7s911/67umAcRLb
KF31g2ZWcB/Skokc6ZC/dI2eEF3Ij59IrB0CNjY7ygIOWy/Yv22lRk7ogk19BGIO
1bMTGMhofZzcDJ/lfgtBrn+qf+NvCkZxSWMDmyev/hwVH/p466lC2WHMerdr211n
poNicoZPdEwFnb7e/3/A9KpG1pO2KInUZHn4r3xQpM5upKXD+cxOhizosx1Oh2Ka
0+mBXO+WaucZbRXf4riEjw0wjbOcMecAmWv7EnnllF3Inz98wPpqTwA/AjvhgtsI
nJAPXPt79kiVJLevDEtHgX1exHcDOQe5s2d6+LC+S2iPylK5ZY/aUwWPHHbkceHM
vkOerKvSRO03qGjK2cWeilue+7aE8170UnmWtnF/FE7oNcDyj3hI0xhN/HyGMQkn
KEZxEF1cCfrv3mefTtD5N5Mi6VRBsTRn6OqWwG1puiRA47PEQmAkqc4L0jhQdM7r
qyHvnp/d780L5y44Vp6HpCMyDSdOlAmj5tnLgvHFqZTQdnKTVUSS/O5AZ4UdrWTF
cVcG+AQvp3+BihqtqSkbY28GhHWwREQeOsBBpU9Y8snx1A0U8hUNC/YnrZ4v0zmU
55+Rg/oSRamc+IE9eV8P0S4ZgbOeGttQTBRCRpLFngGZ+4zLrlHdbYgQYzmI6CTW
DbCK0lGHonL0CJRxOuvXSARopfUGeNaVZsyMF7ECizDR29ABdWPnjweFvL7+Eyep
uiuMPsZUl9XXbc3r+jChBTYSUPcvnU4TKBU+DvzMXxMPFKbJBhbBgreMLK5FBue7
FVETskxGf48JhY15hj29L/wnSgB73YFV1a+ctq30EcWntemY0rbEoO6aIWpCQKdq
CJ8CxBXoavjfC4sW/mQuboR41smCLEFqKv3mJJucZUiXFLDJkWruBz1We8XxGNWc
S/TEhX6rjehbAWzwVFvaNvRSsXfvCa7YePJ70RexRKtTpOmsqVDMCbOr3nL+j4QP
c6mYfWYaIBD1REqQ4wPph86+rHY6sM27MbJn0bsXavFVN+y3IvIeLVvg/SDv0YHw
EHeADs5jJKhDTqo9a566Fj9tPtDyfR0uv2c/r3fA7JaS6yfczGQbVAXGxOGrSLpC
JTUaFve8BioYAjbLKamHCKfYuYHfLk+6n2DwK/27Lii9tL8Rabm6ffMB83NgIdVi
ibUK+CFH9MWd1HMr7Q47sEZk7BBsuXHY5FsHyO1vOPcCEZo6AcBCH7X91ZzxgF4I
KHR6XZ8QpuGnkMKpk+sTC0PRyTtHh3TIXDN411n4pt0DjBcnKLJIIARkc34aRb4w
3hqBbiFvMaBBeoE+j1P5DDpxpk6uja9zhvkQK/umQOwQ2ktgPS7P/TpuO78v+5N3
17aEH2PZhkdI7j71AtI+mVs6uHQUcaI76atbgZPobSp45/yeMwYIFDekbBlzl2f6
2jJdNj0zpcbKQGPSMbRHWGZIYGsXP3m/3dcfl68hJHzSylGDxOWM9thdY3VhE3W/
Rk/KrdROhtwvA3YBYJBYaoQLi7Av7ik37UGFfTbH5w3O5NCzW4/dLRKCI5BiiW0p
gtaPZaBMx/3yDXY1EmS4nEBuagiRw6q/hcaSq5nAXTLyD2gabaeIS6bRiZQMqd4r
XqzFaIPQ2DJdHbd5z48k7zERMlN/q1pDydj2itW76e12REpAVx/+BzT010AZe7iG
3x6Iei4imd43t08Yr8hVWHVKOYLdUE+ADDXzjFNoLp6WS8yc8AqSWofJqP8sqYv+
/zPfyaQ4Yh4T/Wk01EGn5F/pw0Vi19UvMqQPHT225nmsMDbXYLqNt96/pe71QtFO
MVq9eedkKhTsk2Fz/b/tELzdDRxhRORxI/AJGUHwPQL5HnRH/3ClmWZEjOyWWzbS
1AF3zfBCSm0Qf14XtZ0mVTw8y1N6D4P2SNhLlEsOY1Ug8ar90GTh8d7zeU1kgSzq
NbATEx9yGvNT4WfUDTAul/lWszfxgB4I37UM9AXosJG0dbLGOg5k5Woo0hULL1qX
u7iqQ0L0Jupvkgy0InYo16WIYSIzS6zGBliA4BBhlbs95GV/p76aEgvB1YRdOXn7
RDQgumCzEQz22mNbO3OsQCCUioJiVvd0lZd+kB0ZiZPdBriDF5OoebKr5DUGqHax
Rmd/Jr21Ajkz6HkOrUeIKQc3UprPPbXwzZyv6Q8rKTzdgpKvm8A02885giCJvED5
H+nUUI9hXyrxeDyLik+XaS5lj1wT7zr8HKcOb0EIypXuB3QHTCLuVckEJje8Icwv
1VKCFntrIcSNwvMrq1P0iz42AvrMTt/fAEgFGMAlyMqRe2Tb0/eARAJHGdrhFM6C
dzohLegA3dQlg+lOb+mt8zgjJ1e8KdKxV2gGc5xFjncRlRLhKhQ0GJOpJKq40BL5
TiOM/4E5l54GGsjALnjogA==
`pragma protect end_protected
