`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
aihShEwC+YCmtiIp6dyqwlLARnX909RmNFkMW3+FZnqKkaGLKpDuN9m/+5Lv9qLY
P/dO1CXDPd0DSNfW+94i3Wm+UknJpR9cIUhwcQ09MXO+6SBITyDOP4mDt5UUcxte
mczsFe545Vlpb4gTaIKKo4BDsmu3xHnltWHJArO2OFedTOxloHv8En9dt3gFyDg1
JrZSEoRILe9TCY3gYcv8QciMc7u2monShlBgsc2493RWDML3LTrXcztJwigL/1L6
A+klNKkc5EKkRnWxeJXTUJXZ/mlsoPnA2mNT+Hol+zzxHKZOp/N8j4DorHfwvCtf
GGJGkNDt71b9eAMESzJ8QA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2896 )
`pragma protect data_block
2xS0xt012SgoMHSV4VX6kAkgJK+7UX9JgXJmld7wp0i1ntjtHZXyyg2BNLg9WbxT
2syrpA6+pg7L6S5ikJCXcK/GsTLv8m7Neph/qegr4fqICXN5x4tkaRJTmhVuBfpG
hE3NBQFULbIyI0U+7vb3S6/04fF+P/tJdpdZDJKDz3BYsltE1w+7ZAvz+0/rf4nQ
qqPw3H3el72DmTySmQY0TsXE92fiARgmRpRp0QH015mA9fJGF/Opdr+uhuNxdpik
GGh2hSaPW5tH+FgD9B2sfcLTQQaC8/o4RNV9EFOk5/zsFE/e5vBiGkUzR/WgeVXR
LJJXKvR5xwAlZDcrXiTLjYE6k3E9dUnPrCRuaei6MgKOow3cU2pUNGgGDIooS51n
eGVfXB2Jv9vtxiJXY9Kew5A/e0gP1m2Gnv0wn1TG/FQxuAvmS0E9Cg5e8/PtHWKV
jhoZ+VYwdTI9g7a2P/7yoFxMg4xNTIj9XKRk6k2DxyfP4OJbf2kwHu2NPxKT7xrm
9c/Icoimvv9xCeqD5UEEZxyCoVyxHcRmcRa9k5/frKpZA+jFxJtN5OQ+usIXrnIF
wIZBZFfA0SwWCvjNACtwchQNFll9SKF6xKgD6oJMFqQ3KnXhrCO6GbgLY3h7+3Op
BzNIclMZlEKgfMfDsz0icuYrMqLkkbOzklmr4eWPxDxxsiAsXLzjJShwPL5Y/v9d
8V/ljJUyQm/0P0utgDe6mOyA6HMSDHMz9pY5y9hEO8b8N6uV9o9qRqD5UfljTLIX
wR0h8CCjRMSTPuwCAdnmUndD+cBdQ0PdyWNGQujUyOLwH5qqCyUB6w7ZSs2lJsKu
g5I+/253R/pQbzx8Y+Ucn16NyQTgOih1cXa6hjAtK1v749YRjHkkO7yjYyn6Uz+Y
xWdZ16FaaHlWMm0Xo/7cr/Cj9o7FqCWvKb59nHrhBlsXR+qE3SyIQ8svcsYZjXN1
oTKxefVXPNew3MXVNwHRbHlAp72zpJqUoPMvuBiOi3kvum/JnnlsTKosFGDj7GT7
MwD2chGGFirF/t6pCRGyN768FQ+zJ7ufsviGsshJn2UB5JyuNWiE4dhNrwcq7aHn
YDy3bljtJVg4MP4Lf/tpxnqmPraZc+3KtzRkhuIU7HP1T53Dy0gIF13MLXZVeNkq
QyCwO8brTs6Uv2l+5DnwRf7odjX4PagWXdl1e4FpSGXe512YSkqwkEtKsi90tWhf
2x0HmBBxvYcLOtDlV3ARJk7s/26QywH6ecUUU3j8H2r8TRLGbYTc38q/BfP8unX2
fal4Zk28XzXrP4G4C2Y2ViOhkA6+rzivmSDUdayAA2WyEQX+JaGaJhMwJLKELZIt
R6RMqPDKQap0sD71X76/v/bBH96gi8+/d44ChxB4LEaCGsvLp9HJp8Gau3Y+DYG+
NAaRyrCRJc8xhmsfoIMC7moM42TyRZiX7+Rh5HWL0xULRzn7dDYat1ptB4g/D66b
F0peAao1Mwt4fnfucyw15J9Atv8qcAGFmE545lek0n2cblZkkySgqAFqywQ7Cgpp
NeqwUgOOkUDJQ2E+WFIdD20xVc6XLlxJenprbw9ktL5f/2iuNu/rQGZegC7Ip4qh
5gd3LbACtiwuD8zYA64uC+m0GSzp2pcF+8+VYulhNzKP7rTyr4HvsTs47fO1v8y9
xIHaxhK3OkOy6RCbK5uPxBBiCKXbjvGg4BAMXUYWDbXnJ1Rnp2TD/d3fhEy2XnAB
36aa2AH+cWVlJtLnA6e/Zr2/iu5bvPtJPd0ig4a4uOckYFcWzaC1vizn+9Lkdoqz
ODaEenve4xajBicrNXKlW/IW7RW7VdIoA5xaHBp9B39JUTCmjqq6zl0OmHp5zP9k
t+Ni6GRi3BPDE8ce11UoaSTVidvDTVaSkgFXOBZ9zj2/l03dRpQyWW/9gVg/LTjK
TB91/BDjfXtxc1fHsupW/EM/TqY3Kggy4lEvoIGLqQUx/ff77APleXI+qB86/SMo
C+BPAW1ZVRY3J81ckKzoDX1aZJTZfwOBAIKwCWGrxox8P6z2UUS3Mw711AIscKuR
ZvkLia/kwFntD+f2ftcjCsFkBOeEaFTPi57xlFDyKh7Rua1wd/Pw6GLamzJkWmYm
WS/2XbLlNcuUpblhNhNGMyzuBhXaTF58WH6kTld5DozsHzBmgQ+Sgwt+6tZ8+NQZ
LosPmXSZ7PIh2YggPboZhJ4tQRF6CJe5vwxOKvPGKQe7jHnVjvn7t2eyK+8N9u9e
x64gfgo3Gyib3OQTZ5/soxWCndpqEMLU/RwhW72nBu+WW4vqr9xE110zbCI4M7Z0
i5Dox9wMq0rpW0bANR9jAZWCrITU2iF+8l8xQARhtFmZ/+Sb8kD/nbejEY3+JGs+
IDTuRkh+cY87fsU2gal/KTZPw4JopRW/J3V8+GTZ6kVGijSeyVULJHEh76OTzZ8f
ELdmiRr6WwTnvpt2iIGJNDvli/bQX9TcHfnJx7/9FrgSSYHnftbEE4A3r1tGowif
Doz2nxdUezz4KpYZUpbbdi9VllnHzk3EBvl/lTvffd4oEkezIy+G7LqhoPl4Td+S
CWYFSnm09vsKRi5E+QYM4Vhhhs09r6LvE4+dBU4bEU7l/3nBRL6l1tTuKpXonl+7
g4B4aHWPoj1/XYPEV4z+4Rq8SkLuPcUHysWkOsqr2Joz2oAE5UsOEjJmH+eg4QXt
LmTGTGtpRTxjUNVIg0gu20+htBO9AZy3n3cRk+qt8KWm8wAQKdjiDrCpjfDd3OQa
Pf/6mPJE/kD+gTm1UJC62wZtoCHKAeuw6pGSnUhGiFMJxsR0aMRK3jYDqwESf8XI
D+A/cSdQKB0mxf78idE6AZpP0OhUc2sxWS9+LIJKenC1aTjJDCiPNszM6pcZhoMu
3RMkScYoXcYlFfsjhgec8W+k01cx44ayeqApJV9i/CMmkniCnxUJM1Gy2hI1swy8
BxBTx/pR7GVWoC1+g3WtqMmga6Cfabsdv+mYTXefqBFvzS5E2/4M4O/E0/ZN/Hdn
ZJH2Y7v8kvLwrbiikf1yf9LUwUzkw9pvXIPD823EDx0m7giQnz5bn4p/wBawyNtQ
Guq3pDJOLaBJ/qioCvC9y2YaZKWLTZ4Z0gQLPkRPXMCvWtLbkzhrCoZGN9hpXxPT
Twnqcl0yx0j0gwBMFpGWsIm2ofRSybfo571cUYOjCVtKx7DYtSjjbPVUIQGuCHyh
63kQVrWEhyVwJi7347NHTaj9L5DnQvSp1oTayDivmbU6mrN9aDmrcgCiL31pOfTX
kt9qaWttbdlVyuDxyXgga7w4qfKpZqM6hCxNkCcLVeTOxxnv4L8NgolhgxX6HWP6
y2IOetbo4fYrNGBEBiC0cB9jMQiElIDZIzezxi1quF+abYxOhKTpiCIrsuDSrRfg
6g+BYkc1LPQ36APOOFt0q57Bn7VcMeqfUzS5ujHYk2r6SAMkhHJvBaPlGFbeA321
O+Ny665AylUUPsfmmeLO/3fcKA0H65mEjGk0wIa3EfdJmIzpyic5hJmMQq4VdUlj
dcCfoAvUHMJ3TX93IhryLYYtVlaAZNFCXpmOEUsABP/7kFTzS/vnEcHJayxRx3eo
IC1cYphuYsIgFuokHvRqQ72EqruobuPxHGYG0/i+Agy+0RO7ZgeFhQBwtkJW1tF4
b2Nq24B3I6M5e8eKGhD9c/nwoXQZZ08bG5Y0Vs4ks1tSxrqp1OPWhcx3n9EP+G9c
Q+I1gEEdnE6249AE7S+YKTaIB4k/mCRRZlgExfS2GsN6M89WGoyRyNbS3KsAPdka
u5ldgPAZs3L96WBEIyVv4jdThqwYrJ99HdEZQ1rTCnWT2L3EQeun2TGf1ELAcv0j
d7STsN6KnhSfJrbtUxDJIw==
`pragma protect end_protected
