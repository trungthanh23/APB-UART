`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
M2HUyGk5uKC2EPmdG59JWY/tLH29ZIvPKUzzpkFAP4E7AuH47VgxHK6EdahHaL0w
CW0OntpGJXvlfFEVmmwIaIes/nDSqkS91FE75hljNgGC+Q9K5y2X7GJW4l1dQO7z
jySZ02xC0lsNRU0+gxzcdpQxMCsE0zXNjf5W7zpyDLTRwuGjBPt8AkLlOFd9BzmX
WKOFT7P6/sCMxAC+UbEnuAWq16r3kHrtsMis9AkUPh6X0Pbq3IhiMCcgbNOzzsrV
U5BaRy578FqDfe9S5ZS+yaut7FJgaXK6UNxnN8AG82RdzCfFA8uQ875PF5cAiEGV
Y7NuRVkMIisvGpB2Ulso/g==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2048 )
`pragma protect data_block
oIRs5H3U+HPKNFwzx0vhpCm89cmQoAWO4XjY/vnxNjU3EdS3BnBug1yHGG5B2Y0r
MheeYkoW+ZEZaDc5RDedJLppPlRG/J/38dxkYavPNvP81mBSXy37KghYIJHj2l0P
7lTN3YaSwLivG21uTCgzGhF5/+QdLh3wA28sc8S9tLiXORgxM7ka6I7oq6hFUJwF
Ia36Htme0G869LLT/MTVNv889fIIWdZ8DWQWWbJLq8cKkImIKuPx6Htc8Uh50dUE
5kwVG27NouU+4ag/HQbAx2fAWOFOeZvAl2tbkImjQJm06rCy1s3DngY9guWuXuaT
GR6M2eyYOnPDyR2DZ/rW2vTd6E+eIjFAbDoEgvuIWIOWtoGImlh0f7Lja+itdDdc
u+v3QTqNppF3lMYU6HMo/HgWfqPCx4Xyq51ytOUscHAuvfqVjWo7r7/V2V3SgP7J
vbDxscar9BA1wlWfy3Fxe8B/4urH1xIMjS5FR7tkdVsKxZAqPVIAKDfcg6l//NmO
/bYNItNhHEiU5Hflpgg9MIOAY3okHxLH13LBSiLY7wHWhHcSp5OYHWDcRDzv6OFl
lZnkHeT97milYEO8hNlChft0Oi6TdyqVz2nFRQk59+RYpwbSqEK402x/jH/CZag/
Z2YRvsCDC2Hv3GUE87aUI0UAxnZjFv199m7zvSN4Ir+fJr/cEdwgQsiIm6+z/Qsy
aeffhudUQDevzETEcvQSgkHoEy3onRQ0npDQXl1gqr2CivESU1WhQizn+LmmD4ta
rn3I0hmWp7qZHgyKvp6v6e+p8OumnxGEwt3UB/UsqfhhXwG6gf2W/XeN7vaqdlGF
ANprQ9dK4SCngl4X456agOxiGdi+NIeiY5w6ZsMhBEXtKHTvD0COVsdT3RU1ZMst
3pbShgaA/A/+4fpqCbvUCsnw/eOgZJFvUlrOIPJbJnyXYKDUkusjLq8DIa86afgF
IWkgciIyuJShy7vwi09PX5w3Ip/lwr70WLFmV1vvFhKV/ifrpmLo06Y81ejgPK8K
XirSaTfV1ez3lKRUhx+DBROsCuRVfms4nkTanbP39b34EA/1TTghGrvlUBEQ1h+T
9v9rilAScEoTdnQQ3gbRGWlfGh6ZvmhdkLTRtyVGMMomVuSX5p5itDliSGZ0UhaW
48wBddmEZx8Vig+Xod90m0wWToEqxjqXM0B9xqWt/EKkbjYZhpJkg6TPyS1Pm9V/
IA19sMNbC82RKgpJ1BTKKwB49mX8avsHEb9ms5W4lO6naMF5Ezpl+nnk8cvqxUQH
R8LWT2JIRjXQVkbGOwl0qp/lz59xjR+Cs+phrP23aPfpAGnCqxWbhTvKWrRE88BJ
jWrLxpQHXIlITgBIzL0sRYP/g3HUhlkPbftMExZEgVP7cKCHOE2doxJgiTweLiY4
Y5qObkXZTPPruOs0LYNYrKFxUAIHgZtr6aoMdOamQ4Id7I5prRoMQzORRUasD2yj
JNJcZjpGrdWIqFM3stuUWdv7k7X/3WTZSEpzu21SE3s7bZ2AmqvgNQjs4XTslNNo
7yyB49NSFuytM7lhg3y7+UFdrMVhP6f7U6IRaJXkgH3cGE/g7eN00bZH2juvyVxn
SDn0xuWx+uSqD3hr/SRcLM9zMGe3TDazh5qtkgL7Eik1sJU3VdsxAjYqtENV+Ec2
CJ7UO2PHZzoEGin9TjMnwfdFMJG2mUFVd5enHQvlwEaouqtZS33HpXXCqD3hPYod
Ld303j6hI5jMnJRwCgsfhbQo6j0xoqJt07W4zJqetpKUe7O8UlDhu6HZ0G1PQVXn
DkTpj+k0X5sL+EH/hzGWKXQXcjR/ZaiVfZTLwrLncZ8icit49aLTOp8YynSZbNZB
QEBmXgnupkzJFXPwym3hKxdSMXTMmtfVDz9VMBhS30XXZHOvM3HJ9YzUnXM6IB2P
EDpe+CAkUiPVPGe0ENcePM51Gqn6OQt8huylMjIkqrpmVwYodYV3Rp+2Kp9Si7I3
qSnCIBOlLIO+7H80tzuY1IKytKRdztxl4bLf49ZvpYIgqHT1S+d5/j4ZtR2YFQiY
pkaf/YxNXqLWZW3Fv2C5GoWVby9MhJaGWPyZ5I8BWo80tRtVNqwqx9oeLAKdlAPh
mXAKyHxuFRtRqPFTS2NAQjmq5PaJOE/fU4/7kZkk5TFJmoxSRErU3eQ0OCCh/Zal
AW84MVUoeUMWwLCsOWGi7aH2UfXNTvyylxNvOhuAgxBIU7G30AM1FaRjVXck8mbz
WifujJ2rUxiNiIgb2+cfQQTWX8QsoN6+MTFweXzlwBJUN+yE7WOwCgZE8Ml1CNHs
idskoIXtgB4IdSR6/JRBZECnjaMb9a9powFnGRbJA1JECHOEiAYta3HFyjc5jCDN
duCy8rGDHMUEAlAgKpGSIayeIWtl5oVmVvBPhCKDkp5WZav7MWraT8EbTywiG2Kg
HE63TGEykd+I6byyTpryzwA+58U/B4unhTdKaIpMDXe5KXZhLC0rgRxtDLHUV/fX
N1UdKwLmgp39dgDGpGtFlyaxDk1WrYEjOu7IvTHV0ZJzByNQfrOVYFCMY2mCY5sn
/vW7GNhvQpOlrvujYfd39OaoG9Ht/Lp1Fl9iKOsn1JYSH2tF3B8VH8eINXAacoI4
xrmiJJYO0mSqxXdF2JyxfeXypt1y5pzjrVuPFnK8ZpSUP4JLa/snAiBTNnLDvmyO
wL+jh0rZA4Konnn0RIp0J/xjEDhNwlXWCTGCiwG5RNo=
`pragma protect end_protected
