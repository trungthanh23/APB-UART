`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ANoz5NBKyos80CzrfLkoBKaB63hxTwb72d4XRWYhhwUPjfJmRX/PgOGLJSekEmci
zwJhbpTPPaQFc0ZsiNfGYTmbXYllFygdtISxaI3u2QCvSob1+tKGd++rTZxqN4Qy
ECSFwmLDz8Ry22VsZrcwGCjE2PyPsJvEf+AnrpWbBbr+VOEjApTcD/SJJjOjmk/W
VTiL1Q09OFOoDiEb+RLgclRQi2QKXjfCTQQO2tCKyUrv4G3zCs2LxXtFggQQp1im
EPrpwyaeBrOn0gN1D5nyYyQfe7zlDp0XtBjVU0P6Ve6FTJCpF+nVlH/kMe0LT6b4
LkTn6EDg8UXzqz75UNxbgw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1744 )
`pragma protect data_block
7sP8WDdqtF/Ooru/aLxGRdnFKMPOIntqc3Hk8XBpEeRXLEiblhgOJQMOWohdgP0G
+dC/CMd5VRaSe0fDQir2qxG2b1fDK8B/Kqmq/oZixmYAaFE8vi//J9CqVsWIysHT
RLM0CpNQtU63w3a8Hnz4YdzPxAkNUOk79xe4+0x2/gbv3o90kWdSUmD8OQQgtIbj
j8DfqyPcBE2aHqtmZDcKkTHTDC7N2dl2ZU/ui+z6rHHBD2UcGDjuQ1ZtpW90Xug6
t3I+gysBiCTvGS4EAbOR05bQHzwUB9cNETF1IfGw2ErrB/GM/qBW6uayAKagDOqY
0bPruXcSdcFGPzF5KOwTq1qIb4wJYIyZGW6JuRCaWTW5YYHFJrxrKkNTar+GPVaY
fcieMK9bEF8aYa5CaEBOQHl07ieiDGt6UXPydYlG24dPh277NNGrh4l1vTGCeEE4
y1DBwTqXfnEcZK3RooyQJV88T93eqbc7QTs2vrixeNIjBLMTDQF9a9GSRxvC4Nhe
0VE6KRO2SZEu0sVuWsb9fRWyXlZPxKIWz1e+jm9x3Ab/KDuQS/e2g0H9EcZdmm3X
eCQ7Xc32snOt+WY2AuNXT1IiWPtREUJ6Tx8CBZrZY1lWC5cnMkLH6wJaztubdjpR
HVOJYrg6CF0i5to83eIITSlOjNVsjkz5oJTDAW/PZok42NHepqpcmu+mUgMRRUaK
U1oBAle4e/tcYAZVO/NzsbAcrQe5/kM4tVVUbWPXsBdxdTosktbNRaNiaXTzeq4P
f/HtMqkmrwn61bkiw+l8+0XaNtzergGpTOeWsG5z9gFgGptwtIHxztBHgbTnf1CW
FJUdoLPFUN59Lb+7qqCcKzocIXlPSa8sQIh1OCGZiilBIGmYfh6iw1n66QhIh/C4
bPoQtSvx0Uk12OHtWX4NwuK6g3+4TrHDVE6EngQQd1uqDyHFcvFt/qaAmjHdJ5Z0
H7HGvMnUGQM1bFXVN4c90qtdlT5LxoNlEp/NaTxfQOmxP4kEvKbxc7lXOmJ7vzzK
c3uMXl7vju4Y9oLQwiwqDMQ+lncTP5QLgOMG3qnNkSNy/XvAQDIV09ofh9W6vIjo
eB1dYRmIh/IZuQDWWbrPQXKRGzXNf5I/ze+WovnZ709vdIppqKR3xWIiBscQWJ6J
F7a5sTMPG213pTg07u0CGIVvLFe8QkzqETcqjO1wFsQxgdG84o0WpgRa7CX0WYHI
KjLIfE9+eqjhOh6L5oIsxO7UofYPp4NYcLnTrWfVcmVo+wVljMdkO3CW+F8OmU+2
A0NHzKrr9KG62We/bYoYot0a8NlC2FOln3DDm2XYl+b5Qzcr2Mc87+7YJ6ZZR10H
GYb9ncFzLV2Ly3nZpZPnZSu9SHdnz2uTJVdU5tjNNuqHDCKUDlUee/ahLmHjkHXG
qGd0y/MslfTvBICW8DXnd1p47nQGmT4c19Stx9WJcDJCcp7b8IUBbUg1M/iEv6VQ
SOUYG9KWLW2x8RDBiSg4womBJLZ7Es3FEI5POEL6HAZK5nOJjro81RN6jESmLRZ6
kvQtCzDURVO92qgR9X7l3pZczWIJ5tHTtmiCbBcljqYwqjT+wAJcvf1oJZvxMeBS
dmP1rI9ArP06s1D+KHeTu2cYp3ODMZEmDv5T0KrGHoy/1/ppbpSCBr16aWDO4Pnt
WFr7Dan2D3vbrpfqlkyN6GfE6OWCxE7k4BGdI+hIAw723pzuF/lSwBBhmlDb55F0
r5Z8Y6g0huBWlRx28+Ex523bsXn1xMrLg4pnIsUYzQsQq3drtNWjKWRv/swSsQwY
caUEOcFjeMRTDG9rwaahj0QF0dsGZvXs8NHaMNB5g/TnmzN0IVwK7ROlR7po+RmR
cvISKltIYLDY4L7O06Sf4OZC9oQdZg4HV1ZzatrPnSchx8lTxvrXcSpSjh+M2Xng
MKk9cnSUEEDOz3RGdbDC/O6qrcLvyuigUXCkHRWawiFdf2hnKZrBsBKTv6jgDMAb
/Isy3JEei2uyFS8eflXDyuAaoEGJAsN8upKEhEPVdVRHHI1iKk52EfxFfe/MAqRQ
874o2ZnNC2H6AWCuShV39ophNyOYWmsCubrV7rJaOI6Nx595qd1m1VKb2b6tsmdy
oYUDrGwvQztsf4MaCnntj8AQkX5G3+bDzsqbLkvYzs/nIE9GslW1uNkuF4Xjlv5r
MJ2FM2zFiBNzA4zwO0DtIJywrf7r2jh3pNPJuTpfTN6Gyx75njKMyx03gL4zscPD
FKOSfNm9R025ca4OVslHzNzlAhNd6I669UKR4MqUzoZdUEvvDntAhYvCCeZtBmQt
wpJkjkAdjgc8rBSpqb2cGw==
`pragma protect end_protected
