package dti_uart_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "dti_uart_defines.sv"

  `include "dti_uart_configuration.sv"

  `include "dti_uart_tx_transaction.sv"
  `include "dti_uart_tx_driver.sv"
  `include "dti_uart_tx_monitor.sv"
  `include "dti_uart_tx_sequencer.sv"
  `include "dti_uart_tx.sv"

  `include "dti_uart_rx_transaction.sv"
  `include "dti_uart_rx_driver.sv"
  `include "dti_uart_rx_monitor.sv"
  `include "dti_uart_rx_sequencer.sv"
  `include "dti_uart_rx.sv"

endpackage : dti_uart_pkg