`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
agcLD6No8vsyoWomTOOSI7g25gigW25CrZhmORoAllGOm+aYVaCAa6AFGu7pPf6A
j/SWAwh3VpDox8lIk8RTUq1g8nvBU/NeKOpQDJ65nfNCigYazFFAl4lD2iv7ctxf
87gMYSGaoAelG/XvUsDW7UWvqA7D7eByQ9EjfgNrn8XX2O1bRa/PmJffcxPUSvNn
SFw0knh5M9YBQRY677f3ROKQFvanY4gIrOz1YEl4Jt8y3g3eb9ebW/fHgYLL1UYZ
6vk0tZ7/59oT46bTzgNF7Qu4hRK/LlG33UnzlvnOUG//jofaXvqozigTgFNDscY6
mUAOhgAMwlBBwKxZv69OHw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1744 )
`pragma protect data_block
TFBfLUreGwiQNVprOpOKTXku3kelPxCOAMrAx5g6zOQT/DktlQyBjT9gvEsWjBG2
k/QYNKGHY1iFkSUnoTaSqGtc2pDPoGY8bWfHwQsjPm27MXIYWoXrPUjcmvsVhI1C
RKpGrmAek4zC0DH0qFbmzIXxQnT15jihFGN4hJZdSafqfm37DaGlH3RaX8ysRwPx
ZONbmdE7fcQW9aJeeeEixYXXcQHVzfnvNaRw9cTSeK0ct3krLvpCWesQo5Hdny98
bN9x83Wkp/y1y6WGQcf2dkdxdvh4PYPctKEFLb3ibs9x+nrC00d8vxa0BoV0Eb8m
e0kUYJilj5oqy5FyhWLVC/a+co8rDXol51qPPnvsnkEc0xYnzE+ToBpkv1uqCfio
xbM6X8B6x5Ohw1v+BXUaTnwXzinIXphxb1Ark4yK4UteZL2hvp491U0rXuscUdh1
Ol/PaECxKVkMgJ5bcQX4nLvwENbz+/dULB0hfQmQK0gVZgIuLWZ5pBS26zieb3vu
12VCks9gjQShIx9OlM3jfueYVqV6L/Ep32jvnxdLhFtH3XXawBJlAOKqTPTx1J8O
n0skPRxxoYx8WUJzI+rZq5CmiV7chpxKw4hHv8mB2Juy1JuO67YDeqfi0Jqngnas
//gsWuF0xP8yasA0QN8kwHmeryMWo6FD24kMkGxB2rP+3cr6sL60Y39moIFCm7us
ZfoJ0XghUl2iCaaa+Ab/osV4wyslxTRjO7km2VSSHTeZqvuASJwpTIYVeVx3pZM7
BeE+JCAo8lj3RMa5eujXyEjWj4266cHRIoZ64+158/tsQOZIBy+JrnZ8IJ7BlKf7
V7DVFOtE8kbotT2npAvoYTDrQRDWoMa6PcVnJ30FiHoA60Q6hKgW4ZPQpvEtK9Ks
2MXLYPH4m2XjX4q6uqBMTCdaQ9ogAHbqyUcPo3fD4lyZ7+GOTIPclk4sDAhQFKW5
2QsU2X7EEz5KpaXX7AgC7z4A+efET6GiBcdcBSrGorc95PL1HVWPscTZDXETPCDz
xbcbovJVu4sm5/Oz6XD6DlFj+hkukz/ahkOTPGuwTGRfXX2k9EMjk4nsnk1al0dR
SozB/C7NJTgup7xgVat3Kk1W8r2fcCk7csxW/F4SRSKlXHXxWjT7qqkgVXdssE5z
u/grHXH4XQXg28wIB3N1Dio0FM5kRRL9BqNZnp970nhCxn32cAP0ItG8pSJeEFSn
6M8/fFIIyJ75uSsA2ekPwiHLuR36W5eoEE2LVlpMwuYmpsUDvUamici4r84zzTqg
xPxqYN7J0mvjB9TKdxyxmDQeIYiXdNovNRzmNhvhdiq3MLLsSdY2V0efOnEIpVVL
xqBOA2evqWA2sSeMzzy3m1rAsclN//zLF3YZ8Aj39map73aJtQ5QQG0yVan8Ev2m
Y5ktE5q2jgqCqaUk+g/RmzuFlfox4ruKATk+YgLl+pV6DwzUgFqSzWxkcC4u1/RN
BL4XWmcvf4h/nOG+EAaSvxxgpxKhBNOXFmERkeemc/MmxMC/LtEzm9k2etUU7MvY
JWTqoTbEoBWNUJ3QE82P/crhf1WWq7fPLJjy1nm1ciBGZuUd75hT125lovy3oCST
aagFJtKgGUx8wwjzTPtMvgf7hMkqLnKmGjYqZyHhfgt6enEasryMRZeuZI56GvUg
3wQNZQpmtkPQ8VJ3Z2oapHXpJ5vHmbkbfzaNGf0IO0BRKJ33QeBUqdxSWwQGG4w4
329cXh93ejJQQpGYpBC36QjY3+mMFh1USbtJzLBPNjxcOcdvfH+CQxOhdvRzxpQb
qdzA8X6C+HfIhTOvdX/R3+KtSE4ItprPvb5rpCsSvJMtKMbuV9nvLB80xDNRvvvJ
7joKqDMdxJb3FmnEaLZzyrZJuDxJiMNb/359ALOd3sgU3qawPVrmcdA5iN/ahhV4
t8g+V4xf2JDrvXQRBIRzwp24Ow6NbpSG7ig8/PXfeGiQ9WIlpJv1VolMBvI69jjy
B/G5NAIo3ypAvh9p8p0bsKeNEQ99wsPjof8HybIk19Vg2rkHhyiD+L5sxCQDwUaJ
B/+yI4bB8li/DjIDpi1VNNBI9gIep9vWi2jVrJraw66qr5dGSzsKxpXYeflVXM/a
bLa9rhuNqxJO3gzerJJDMEhwns1nFN4CJoaRK0JpP5QuznQAbji475jx6DxXgLNE
GhifWkthjqULw+YrUVaEArejj0sD9oAMPq4vTvK/9djyH+d95YQCGNGa4TjdT59B
ymq6c17Xa8gT4R+PNOjoMy7Zni5N7a8nodH/PT2mUspDHwzowq+h6RqSAYR7A218
PFGvycUHWkdeFrzgAXwVEw==
`pragma protect end_protected
