`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
V1LKo28+a6dicykqqRHuLfxz6pUEzKnvPbjIsb/fW5T0u4e+KU/ohoqeAqC4o3zG
mritYA+KwIiPg5kEce8MGidBAjQnXDxfyGtJwT/rurfo8iL/LQ4VWG7IGCF1WiuL
off/V5LenI+C+Mcyqf9z410qsUS0HvRl9gZ39VeAtRyIu9GG5ihetHvHBtz7E4OT
DO4STkilkIguMhVpLkMtnotIXPxBZKkF+/ZqsToi8jb/qnxqPYq5q80iwdIYnj2W
XNJzGh8eWiopiv4R+nfEziYqZgp3b+bucL02YBmpn1EjCGrrSn3UlK35NaBB4FlT
xbII7WOK8leOc5KPRRV52w==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
DyrgtHeG2rbUuVeOVJ+CU9ZGPHxvxc9q6ATns2IMqmrA/mUzsfXEAXpSTedAG23N
yYexQ0E/YIIRTvni/i02JbZS5v4vc9fUoSs6pOOlb//d600D/NarP5hLdKJlLDke
1CLUE+KKHFLkE/U8uV/JYcQfP+YtlVIsd2AdjjJBySI2LBbJxeLFKeQOY0oMzUYu
YAYnyXYBZsfFbCL8/VXz4xFQjtorXHHgrTCbkaTHQYgO5qohXQuTgC8apJ5owMLr
/QItTXg0zw8dt50CqyZY7BJ4qZe9dJl5EvPAzDi7HrAlWZkdR0BF8IlJWoBWXPAc
1kPnvjYVIPWStWM/oKtDyxvWDWrdhh4vF8VnXiMpvIFyMXO/QbCIY20W3zzsMhkt
p+eOldMY6xBhpTIYol9jPJUjv9hcSNpCo3OhtUZeI+AnWtl5Ex0JaMnbL7R8Z2nR
q+0Xpu88vB4k8YP+4pZU6jjSK6OdGvy0RU5oaUvtaH3ZF+pguS2bvppjNi7oReH7
CKTKzC9yGMpYqZ+RCuPPe/mi9uHG1ZdpkeiQnrRCxGI1EkqohifKyFLh7ARP0MUf
KdGbaxKHjQhvV8j+MCUqpfPJqzvFznmdAmhPiTcvUopsp7qSx7GurIH2J9kF+KGQ
6COI8Wx+byEzswCOvLIYF9Or7REJ1ZwO7eqjPd4GUia7FE/W63d4eDD0fTuhRA/k
bpiTCe5d/uqp30L830mCFXQ8tQ79IFA5CrEgbHCKJyI1rk7ywABV/HfuWZYqrgeK
hGAV6TEz8ssT4aLPrAxhoetjQruUctuB+FVn+mV1EYYNRl1uJJLZ6TvRevdgE8Su
U3Y5ODxHsXYdlaBHv/YXUt/LD7aeCjOB55SnYA5rK8EH1OAdWZ7mgjfRImvUaOv1
L/ZWaott9b39uwbbQibexho1hnXin1dPXAgcCCgJafWOZ3IwM972GSdN/X9b+wMP
qdHRduQr2H1nl4n8jjhEspTGEoRdKvEtNqwnDId6KadEmKlPndHLSYnr/BfDfxOI
E2HS32rnaZhLa5sSJAJVTV7B/TbkjiuFn07L5OcIiaS6WjPF9zm890TS8pTs+tBg
QlygKwIfbOD2YjJAv8ddPSHnGj/LJi61TxoCZoDgi9Zh9wnwNwZ5w8aWRArmuFPZ
sQZAGPdHEdbdm/XxhMVoSb7CsWAFGWK0YRzttbjTIDCczABrR6ib65qq57uybh1w
AttDcZooXMEFftRPXMnG2O7aMEMvQp4sHch+5dIogcl0vNM4/XOmZvuav5b5YkXQ
YvxLfPsGFCR8vIxuKXacHFUBHa3k4NUyVlYi5YCud/DL1QYuwosMMjIxu4b72sUQ
bxKqamOoHyVNzCTxku0W94g2oKik4/lyoHDjVj7Ld/o2C6XR5ZpTCNBTopUxtrT+
xt6nX9TmLT8s/Vt88f2qpjszp3AS/53LLoUk0KJe7MyEgTy2k2Cm2Upvjh2PAYW/
TlVQMy03ROSREfzFGYBkfgbqSrN/RKSm6VZ053UrmAX1+iZo6dttzm0QmHt+ePee
DrGYl05NMlAZzSJ9dLZHTA8ElrnXz0F449xt9ZUkwgTLj4xM+fERwK7lh1hkX5qP
EcM7eItxHCw++7wiDqKUIiablDHojQ5GN1l6GtXqyH9ZQK4nV2F+XqcZb1JSk11o
CXlPAShcd8MelcyEjQThat7LcgoYJz8+0GX62C2j2+r8Fbhc5/zRYSYiSPozmC65
JohAbNauAylNcTWw/3gAZjPCVGDWkqjqoF42EhuB2fHxtJ2yjuYdgjPX7Ew494Nz
kmnlO7BtU39VYiXmNaSmmBJ0QHzaEKTAYaY4Mj4jDAXSX+3v0qSSa2J5juQRMkjG
cG7RLhVxM3LPFqoaLf+i41zT401VzZreNT2GhFX0sU2Vs9dFYUCCfEAKE9roCeTH
NtFN2F7e47yK7KmFfvjRPngTRL6GTHBaDRjxHszmy7RF4DDOfOwxI2Lkh91ULZIn
sGCNqRjWmjcUdOM76ufebRumlwGFV7c7aWhgMTYGZ+kKlET1asoeY3xtH4MO3e2H
LuWQ40gv1i0cqHxsMhwwZblSk334aRp06/cTEUi9jDqWBAxIopK4/9vlyP7Y6PJY
h6Fsyxs9tHXZCSVyMoGCvF5sYNX+NGNh4rAQKPTlIEuEOixpAGO9xc6Ah4uph64l
M+pRg1t8Y2Nvf50u5CLFvpVgdSer7t0QWWudPQ3xPuqKU9h6mF98tdL3OdeDkxQL
Z4dP92WKVY7TjoBNhQAY1/g0UIIK22jHUWhkl/LBIxf4ltoWg+peIa5gj6pfaRbk
hVIffg3OsqN/CiJea4mh3SmABnhB+4OKX52vZkKg9ZhyYNh+CghYSC4RZL11nrDR
+Zc5uSvthV4oeBP+eVa/+ROSjhXTAk5d6+iSsyoXLFmh+apLGlqEpAdZiLrmlznu
A5OIsqZufSKptKDexqszOsg/lnb2444bxSpft80yrxQu7VYrfwEjRYDiAMvrRtx0
NkyFSMTPO7B5QbRJ32T/8AoW8AkTYP9B/KBQm+k070rPCvA408cq0vV7FL/EfX7l
ZpBgtdl744I5DebwssvISpU7rcxEYJPtg8IAt9meSwDIkrwhvaLWyKEGzH5c1/7l
n0I0Lz7FR7diGEfZoMvlbFqeaDT7rp9cky7FePACgIrbgRVijX+YEuFHiCLzYKMt
eNw4bWTDG4+VsmOFRQ56f+KqV4/vl3Jk3iuHsTDyN9gxf0xB9EQ1GA2wiM5S2knm
bWeQxJOy8oikH1RDcm8VqsG/P3ojKOlYi/HO1llrs15kjlO3MSF6Ll4y0rlnSk8K
dy0SuwRRWOVrghjDgsOWofbcMbSsdrX70C9hfsJmKax4KnmtgYOIF1Cnd/MuJNxq
7zKDi7YqO6wq7if71aETc0pUpeKyOiVvpT971pGZIci3vqQJWP7Ool37D92FQGt3
46/kzUmx779syr2CLuoVbL4mM6ruv6V5PeUa2cR3q7669rTnEvvltFeaiTeNi6RO
ymUxiFX+lKCBxTkJ1VwZ4aR9FaNHBhtO427Cig7e7I/tPqu9YgFkY0SpB9ndtiZj
shbu/uiMT3L7P1HTKt1EhYl2dKGfADtyUQAn9xkgtvkd5EDpo9OQvFFrsoxlNy1l
GeT4qviC6cNLlKfhoAi/hmqKH7tPAqOShP5duURpyKqhPrGsaG/VChNlWUHALBTq
4x7yPnFBTvEGhCHUuoqIPP+d/v6a3SrdSaV7YJm+f6Zh8awt3SXAeZdZ3jxIXSue
PJaNUyULCOxaUd46LplF1SVakEowoT5D81gosRECkY6s8US7Z35vGL+bUuG7VD5r
7OYTPjN4dXhLhiAe8Jwm4yiaTlS26PS6TH3ggcTuCryJUxdmqdGKEvfA6CkgCvbm
iWbqZ0wITsgPNXQk+ORmmwrta1CdBLkExKxrVEWceNSkO2cRF62MZQTj9y0yiTnN
5WOxEeJzvmDSbTB2UMhlTPkB8UfZRzuOT8lZpV3h42A=
`pragma protect end_protected
