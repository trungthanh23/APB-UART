`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jSjU4rVL47f3RX2YgozZe4++suq0Ax6lOXl1PONARFmY+FiWeBgGI75HOLt2sWnm
6l2hm+hrTIxXkhIPPWdAs4kNWTKwnlVBdO/PgB70ADikU1mfQJ78+K9gMz6Eq3WA
J7vxJf3nADbQff15qpzz4hjuOyE7U7d5lprnteOewokekZxH5ji+QOCbP/CgeGkX
FaGU2JpXZZBf5QEzJYob3xC6vmsdDYSy1yh5G/fiZLkxB9POpTGUBiJE8/ztcjzs
xHW8t9WtXNmRi1qYYcZnfcrKXu+CL5TNNa06z7qzDUXirlGMGdaqxFSjPR86VUL7
h/6q5qZtwoTpvHKncaSClQ==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2880 )
`pragma protect data_block
FL1gJGgSyYVftm8rpuWY5ReAilq3FtnYstorcGwOTxHiYp0A0siR85oAP1gkXdSA
3hMpfpyeF9AvGEZYBO834DBjoQvZKWC572LUwGi3s2PdEbeXOo99E73s+1Lgtw2Z
goUQP22xIUx231lxm+mRT9owC4UpdCmto5evw5xd/ScjH43VOHz1jkBdcgf+wbZl
AZ7/Fz/YTh93ACp49gqqjsz/1aylF68EuNvT8HCLeZFUmCQIwGsg5fQreZBqd1Dx
DacIHsgYU7HEpo/Lyf34P92K2uJ1EW3ZPQof9fJ8dCJ2Zb6q7W32HfTqkJBQx/S8
DnD9GkJfCuP5b7PywFj5TshqJBh8/9i732Mz5OdNb+qCjqHkVTsTLSCSH7vnUUgC
EyfYdAr0DariVh3rliLcXCnBHTXkLhwEhGz/9wkE8M4G43sTvWKLErG/Cv5vmogg
tVWrV3zmvYMiOTN+fB21CbOMpmkI6BxpRWL1ebXa/Xz4Gd7lMTog3Va1k3nVDn2N
VzkdjijZVNF/0YAMRjWe8hxcIA8Z0ylonWnKNxqdlwS+aD6DwtuVbpDTH40PLrQs
Z/2f25gmdXLAQLb4L41sNveCFxW/9d9ffzD9ZmnzvK5tdeOJG4DrWb/2MVagprGP
TDT16X3Ks302uPGTKHwslEGy79Fr7w/cvAi9wX87yX7kOkVpsinKOvW+qUoyVkAT
TV9av2DqGEnMZorwgFjXU3Dvn0M1mzcg+jayUZwQA7brvYNBHOPzO2F4/6qKhemM
XV6ySu1VEFxx8d3nNcPLi+2LMLUBrCctx2ZayNR0GvyrPufydkp5OPLUWp07GL9R
rTkoIA4HVR+BJHlSQj2NbYgV8fTzVcf+qVN/1qokYDiwIApCyGOnTDPdMkfxrGJv
eRkr3GphQT+f+CH/9RPjz8n5vmoCc5FnnaKlR/tTc3nXhXsQ2ChsFScl3+lBokQl
YIyNp+1+EBpcaYqcyXo0gofr1rcReNfS3cwNuzRyVlyqJD/mmsyptqw6eS1KL72w
pZ6ErBU7baYKbN+sSjCjSs2PbONYLbdCh2fdycW6s/fN5ycfvkcNp6YGN7nEfG4Q
W8G+Ane5Wj0Lxa8LV+ebUwtwf/02wr7tV/6kriDDyxUfkin/Fnwf31uD+LKcJf8z
OUBhPdd5JtW4XIIkjEsse17QNTV0jkybprEGlTpTY455Z3JW/QLz6KgWdG/KShJz
CogQgVJF83Gu86l5ur/GdTD8EeFmIX9+AzV2tn1efn7ovQKDyriXkCHhQ+GXAQS7
lx+cOqp5PNoxZpCyET7G6siu8Y0YoZ8DRkCKEx+bsofvUJ0JyPblGpVM2GpWCclG
ANUpZTUSEDLEnT00Rl71NuJK1p+jYRU3EEdxzAZFZ7EzS+q+Jd6+bhR+um0oa3IE
1iF8Y1fE6N2UZNPoaoPS7ue5E/Q681sOJN4czsNg+K8EwX6lqNCkyiQN+HHoGUqv
ZU69dj2JX5/dJmX9zCi/hCv2idoO4z2GlqqaYAwNk8UsW8Q0ilZiWis9NMgyZrfT
GpfZbogetPLvmdcSkBOQDe/jsx02CG4VTyjTU/CrHYe9o8GnJ3lNAnlWBq/rnfRm
7n3G3qZKv6ALL0ngXZkx4AHBeZ+f6crM83zrZQT8psDBvBN5XeYmgcGD3ThBP+W5
Ig8vcHNkMbvqjVkV3X7dLMDsZwmEG6/tBBb4VbpeGDHBgjqgtFa4Z+KDoHZJDbtl
kD5QRJaFPimflvWrU2zOX9MpF3iFiPWOOe0JYuk2TXSJmdyVKnzNG58LAcbXuWjh
eefWn2JUwHV5VHuWrP6LrZfZl4OPro0U/Umi/wnu3WpEYvTfThRV98JyUdGQN/lF
x5sNhPfM/HB4fRDnU5riecUEj6RPHKB8ORfM3KGTcXyW7LcHOTIX663IFPMfSWwl
pAyBA651K886vZQEQ2cB+CmrP08dKgroL/S4uUeFUG4ywk83vSfLodYkC21cIhze
E1GtUG9gMtPlbFVDq5B9HhLmy5FpWDM9I+q4yhZ2rp8lH73F052WId+PYFx9ajyD
XeMzskLMfRZg6fsxHqp/rBzXPE2qNHqh/Sa827o6usIWyTuTUuDZGb5s4OJLTBUE
tg5DBw/wHacKj8QAif9Q17A0c8WgpsO03Gkn5hxAYVl3xNy/TB2pV0ST2oSvWX40
MlKDecpuFy7g0XpUdXBXbVJ8FbHN5+IJS65KxUhJop/VwlLYXlDwm+mTs+1ySQfy
CRf3fDhkpVbeVW9cwZQFOKmfHnCxG1Vu980cTVX7kAbc0Zk3XGIAEfuuac/e66M1
3jDR0dO4iw1ffpuaOKz5UutVFDqX5GLzlqyur4wBW8/k997BLjXJ+/IZr9GG7DuB
e5arWEFWR8r0BxELlLNiZ8BmL0ksqDBnBFFbJ3OMGak7mVrkS4SeYOG4qQEbOch6
sGYko5LSzWlpAUE0EQUv2Hwt9fSniLjGtJq1JkW2npc/JUiLGvwEb/crfb13bvNx
bUEoFb1aYtvfuypQnqdNX1AoIg5X74KTRSwgsKKxy+zzGWK0eaYz4Br0/t+zYlxy
M5/Gs0vBzQocyeR+VQ0BqlEsndGW8f40s25/Vttv9IfU+3ziiL3aCGEEq7Whlot9
6VDvqix5zS2oAjXtOG5bL995yH7vZaRZK/JHjq5KBCpfw1HhUPf1DdhDNIn5zV0d
J3mjv+LQhVCOXCYad4gETFlacWLvKdnMHAyJw4psFp8k6u0YD0fi1pycCRNVG1pk
vBlx+4wyQJDZwWsXli/noLHf8jpwaceif4fhzHJsCLG8r3WjqWzsO+enwFwhXIC3
cU17yXb/tf/LZfd+3e+pX4sVy8n5e+wG2edCBHG0ZlpVsX6hm8LZNFVNO1E2Mj5i
leCozIgKH4XBNAUpSqotmgGJqjARuZ3CvrKqGvKF80dUHbEkK7LJszfgGDPe/IqW
HxW08XCIT9IUOzLXYWGkdX3o1U4Um2AOkLRNpBT/lqK6gMPXsAmGX7KEsyXK0fNk
EANwAadfV7+sKYDctypAtvZ8fSsqSUHpWgOq0JpZyuzTO+3VrH27QKbyYjjo7oiy
0x5Ap8rltue7/R/xtTgALTkgbO1kq1/uLcHzp2TzdIPVbRUn1RTeCefFShe+W9fj
IC0gFn0OnYavcanQw5eRieRt/UZhgpcPLvys0j43oWdhIwbhhh7VilXDUicPwgw1
b4x2cyW7fnD1+NrkIIampGxJ2er0f52y9GG+xTBKijFfprspP7rZ4K2BFRaFAWkW
mOoAnRazt6wIwLc+PGNIKMVWm9E6W0J0hGcXHSeKW89t4GWRvVcrk1PWDQJvVo3n
Evop8Eg44kv/zribpAfZa4TA14+fOZRQzbdvDAerBzPTS1gjRw86CblE/0WHQORA
pA7zL+ekEVQsqs2CHn8IUOC/CP/vBcV8vVQNPcC5+99auJfdX/4F4qRcj8y6txiy
oUCLib4Li0nxObH07LTU0TBABpp0xixohdV2ZhT5eAppJ6uxEb8E5va2aM1OVJyn
kpuI+v88YOpnJiRihczXq/O/y74lDpr6KN1uDyWqX4NnFt+wnnHi6HY9Z0c60Tn+
hCJoZBxgz+vatY0vkEmiicttwZ4v1O6RzshocKfhSW7vR4hqgsstcaPyfF1a2jha
qzro4IrjgX5OAQo78MBDBIxLr62aQKy5ANaTFGv1TaYOkT2gEIpQw3rlNSgIhEsf
QMTdYJVRIgU4j1jReuaUPulnVvvtzV+rPn1XGdHFdSgfaO5gP1iolUKfNFb86y+Q
cplIrP02K6B8uKd5YGUUZUj8U3EsPz12dOHmEZ/w7MhwQRQXBu4oA1WpQxd5K9Pc
`pragma protect end_protected
