`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IT3tlgzruRtbAsZLgfLIDEdpICJ/dNf97Yppsgv9fJbFiOzl3t95A5jr/MuwCiZf
4tJ8rmdEjE3ummDWl/egHEmFbtpbrWXjEfkeCsCbofRZgEVsAaDc4fgtnQ5V9GL4
S0pD5nmXNaJ65ht+r5UeWdbofTkFGgre1MHcaL6cDcNy5SFTwaIuN6tZrpFuTKIr
eRY0cMlYRjCZXXMuIYena54tT91R8wZSjswzgOEpk5CQ3VfU/WrEPOsb9Y/MfK4b
oxM64+rLeoubNiIUJerK3dBlCwKM22z6m+W3UjSjO7UnXMH2BvUMcEf/O/tEcHbi
XEGoZacEAkqoPDjMhpfC/Q==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2592 )
`pragma protect data_block
s1ZFBdSq9ksIjqp2uRmOdt0lDEEAvKqf5LTLNekExMjDeujBl4Kgapcjq5D8ZSwu
CQJLkgJ6XZOezfSWSS4pCkHPCkGivOZAeieoNZFdG9TjDBlU0iy2l7sbT1LjROmZ
imId5qia5breEaoHA8V9M/nqhpBbWhLw2ITcd95eCkQcwClGZZs0AEHy7SiovgTb
1Z3Sl2Z/84XKnlHynRo5QNw7Chj8ybOpfK8Wp0Wg4vgOaTi9ttIthR4CbIRlzdCO
GHS86P9Bf8WaSRY6e8NO9o8ou1G+4RoZ3PpDVt7/CoS+MDpcgZBTRgsbYir+Wk4D
E5J8tKnOiEUn/2Cmy/uTp5ThRtQdhHgYpNIo8wSGmrWqtwcR/JGCAoCAMQUb3EEC
lfaHa9E3DEFd/FUL6xF1fo1RJysYJIkPA84tHOMjqtzVSrb8mfm3cdueJZ0gUkg4
8fuKjzBsFFmRWvj/YZfxyKZ2eHr5u7UP4DLFkDkcDlYWPjhphjMBp0n9vNZUpbAp
WfBGPBj4xDmXxLQyGV7gbxIyYUFLLH9g+aDCqyyWBON5W7CUKgmBSKaC1wBK4eCV
dFMVL5N9cH+XOCebupvZnJqeG7WjF4Fj3WCVvJcE1BBO/cGCz5+anW1GyOA70b8B
4I+AqAImRVaTz+1ijwbZUY/qhTbrEVq9wByVKp7Kzp5rGOksc9QN+diQM/7RJKkw
JlX2NYa48GqaBICNDzXP8ZWTcxccqwdsgOPXnivS/RxLzfHKwKZtKi3zPQYgYbaZ
+J0YHmrLkgU6AfILYhjJqvK0fH0qalcDznZGtxMUJebY0uCcA53virZLvPvmz1Fo
Xky+vzRoX8517MEa2g5Ctz/a9pZ3wq/laXuBSb+rZkCAGgIDVDccG51ogktg6qO4
4U6KSMmYpTqJcBN3T+A2z94PTVhqk8I1qZBKhQxjMCFDEjz++jccDW5kg6GGhI3X
N5Bi5AqipMAGLPXaE3Q6lCAxHnFB7wfGsFgNa6jik4dZvW+OOLTFq1tfdMOyHed0
uy47SDajh5Ou6zkXQ36uPzhZdSdOorws4J1V0Vo8s53A7x9DptfNm2DuHu+LcIEx
ZsV3ahVbD7BeQ7zEyC+jBfr/WWHRA7o9miS7qfyYo5h9oJWdUKz4GH0AeLEAJh4H
RfHhlRis+TRY6CU7oGKjghIM+Da4OxtXGtRuHTR4ICY2vY62iXhI/RpCUVqrmmjq
9cwjDzXnRXGW3oM9Hn9I9f7qOb4AuDGjqNI2WWdrU/ursUbgruquXwnQB3PQnivh
HTt63b5pQ0vKIEIZ9FfTyR5HgCERUCySAAYCZRsFenJZA93UQmcOIfGw8cUXjUhW
bPn/tBRMaFe/0xCZFCDnuPBff11w5/uAzhxW9ngTTY1wp3XOTCAXrAKhC+lOF84f
B9FLO2XMcC0eJB7Tfc721UK2JN07KlgEomeQsRuceQ6/4Zm5GLM7z2lhagULEhrq
sCEDQfXYlxAxmXSBmxxg3ZHs2jdANl1xWdk6yNjMriENy15+3+uYbpP/jz/Iv17g
rlWnOaEgWP9ubkkQH37/OCQnustj28WtvN+/8aEjQPCYnr8HHjmaYoZf9SHqQgJI
2BN3CLtHn2bSnJveR1GeT2WgXp+MSyq88ViqQXsnj9DLR3QfR+pGC/TbABx+y+3e
WCvOgIqEB5Fn6YgveYXeil7xh5//cxykqRZdtBPoA7DVb7fMduoz3RTdKkxxVm7Y
IklUF5bPMWRwsrOoz4ZUZH97LlsN8GGCSpQ5n63c1fVLU/E2ww2YeLuhXvCW8GXj
5/8xMkYUEs3kk7O19pXaMBJKxZgZ+ZG4D1F5timh/Hs+wh9RD/9gnNN9C0qDBlvQ
HyRl08jaDrfzfrepZjSQ7j8zY+frTWWaVwiikc931/FcbkdF3lEykzxWd7bG+CjW
FR5nHIvl8wWXfRQIBpuUU61lX7kcuHcPO/d2NvdyIrJHAPzJGycaFdiif0aXRllK
iPcRnkYaKVOrDJbbz6BWDIF30t4VnSSHEOdj2ZXacSD1XDvMi3dAXA1nfKwCA1xp
kJcUAoAVFjweqYpVQ270rjfBdajmnEKb9W/2EScvj+wUcTcNrZxuyylLik1dFp0a
kWNMrcsRwuvuGbz7dJ1m2K7yRIja2HTpXUavVz8fRj7M3sdUZrYHydn26Qxx+dzE
8sw2NGHcm+qwQmWZ+IwZpUW5nAU4ijcw7RldtRkgQoE58NzbD+p1AARQy66q9W4P
gMGO9+RDb8ts+y90e1HQBRG9y3A8HjwNmek9ywMqAZ9NBy4PLoF+WSig1RJMiPPj
Nf7+W3J/HmO761GF5YWAiL1BTSNEhiCz2Lq4BMx5smr/CkEqta/ublaVX+WQOEib
pFfSOZoGXEY0Yv+OnIcmRwvKi8iKM3FPTPKf6ja/rmyKSc5rSc1M6HpXVcrpTMcR
9OEo/HJc9m3ySzMCI0rjLLKur8YOWSrvJlHSoU3CSaHH0A7y4mfjgmWfdlYWmfvL
bLN/YkurZ77nzxY0JV4jwZw5TrrHCvpIk9eYaiqRa4tqepehqeNqKf5FZEFJ8ksA
tPSeSK5OEuTSbZot9KjWXoD4iPRSfQRP423rliDSvhC/drSv2n7wwkfeIODbZhzu
1O59gB0rJtpv9uFSuD1mSABQ2fIZu8djLihzF0X73UEbygjmp0BlGl4oLqTgfGJh
4RnQ7CwRlap6PjBpkltiif/D1iYn8GZDzygvNvbJCYeR3MOdPfKeYwAwkgcNqVIU
FJJDMmPKboq5df+To+U+GpjWUIU1owDIzemlCmuXFSc4owD1UEaSSOX/bW7DL9Y3
2y+7bIK2d+ZOajUUA6g9jxu1xusIpDFr3zKRh+5WxqWKSEyUmFFEls8naqIc0unE
Zb7Nf6L06LwKMaQFX1QWsml5iqZFlRADJR62t4RJEZzHzFeslSh0ZIrWvHcDzmwW
i5XrpXAKzODgS7YCIxjKAYLxo7/HQXdq2SQPkW+dd6WYueftOCSIY5QaZO5Ehvqo
AKYlIsP0PvHky21mcT6SnuTb+7iABed5MqfjBP8aaKLNR3QBGf1VBx8l1wY2ofz9
8yVdUJQMl8JJLf2mE31qFi5p1VOVB2M0iR7dAhqsm/jtfpY6UrCYqq3hzRxS2TVx
F2kNIj+NIvChzCeQeaPU46pAIssQicEUAvdr8cwdKBVH4QnNgrlG73WmW5MLatFx
fZdakwwwIlJiem8GHEpMJmQ0leJ1SH0vXSMCNaT57KRLDlFCG8zYJqOEyokwhlt3
fRPh2/8bf+b3wXu2Na7jMCek36CImRwqwjg8Bt79mcLWUklVhoeV2IROUJC0+cFs
88eQELXsxdQQrhzx5TNcz+d1tX1PuPYTmbaQjV5d33FowriXETaQKBrwmKcNyo6J
rm8zfrhYoNPMmwu8iThTAWw/AEitgi7jOyhkXCzjtioWxEpQyIB4vLJxr4CU5Gd4
`pragma protect end_protected
