`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LyUMmV6JywTmsC7sQ6qevG4FlzzBggL3XZz7QNLicprpicq9OvY+y3kG63YY+pPj
3LkOcrshfDOrqPnCRxNJWxTSarrisE9g3KP/jyX0QysclNVQ7J3EedfBPDaubD8b
abZZL4sT8cOo7dL95JrisP1v2iZjY7Ms+D+NII25Vt98xDOZpTraDZ8Ie1taxG3E
WC4INYIYI97h5E5v1z0JQTelRxhquUk9XP2QwKuVpY6Pow1kVYc/PmrCrGoMjUXe
B+ZTV06rSKvdHhI8G7CnCpzH4TY2HpoZtWBQoVHBlOY4mT/rzKRmRICeAyHBXhcf
CDvgZi1l/ECiSuJ2Hquh3w==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1680 )
`pragma protect data_block
5/iUzgxFGcWXg0jd1dZ2mX5zBGo6Cp3MThV1UpGpuIec2Dv+1gAWWxeBk4SDzie9
o10G+jked4d3yz7OtO5TusgWaF6HwkcWttNFS4g6cT/eR71GlDHk2+1p1D04Ul7W
vP0eajaFc1jl3Et9pJxExDsMRYcuOscEUNR14Oxz+FlyAxcBNXXe15kEn8c7RnZh
Mbmd2KIFP4Asc0JUwangIqZ1HlxuRIS0cXKOESN2dtZi5D04aFxkN4+hcYrcSXn5
87sbuDbgj9cS9HaPVmFG4Z7vgJ4U2dtktQnUSg0HzXkmNbilBGQi4UdYzdJvLxOr
36zb5dIM19UvNHz+s5m2jETakeq7T0BPd9WLN5TP0m370KZIhiKO98l7Hv/afdhh
QtUU36K/+j/bFrjtrQQ3D59CguIkyFHqoIdqdeaxhWxxpZ1vWLT8c1rFrjlvmitP
aZnesQSzG6yWkaXV1hwSMI7PvHn9KK61xrdrEHoPo6Vj5+b3HDyNCwRIy+Q92bVy
Zsh0x+zkS8ey6jkPJXFLDWGaXxGgwPGmHieA0sm7tTjAhfruzu4GaTyaLXNpsT9P
X1NWtad7MWmuL8cu9vV+FLpEVS5IvdPI59zRKTmvq6R0DJF6Xk+sVUoi8vQOasBe
hg7a696YrWLjQUhxXyBKgMAcxBNLYQtbG1u3F+GnxG+p35TxyWo5WNCi3uXaoJYT
F1l0Omqp2pffuqzChEh4OKjpuPos1oHrQaboj+zZX8w/lr3ZvU0/dGveMLrCuZwB
C/6zl3XEZJ/02KS0EQYxZEfD+biE0KW3b7ru2GS8gSOq9o09/Mxlad8wJlfMBRAY
QX2BvoiBGWBhLZJlRvOb+PZpjY7qbrqFqc7vZhHNaLIdKhf3mmqxhwGnn/NeYWri
Ch+ZD+9WykC9fibq4IFC7VEZ+2rTPvEIB4cBTnyh3/Go9AMU9i2Bk2gOlmxXpTz9
aupKKjHHgIDO5EmBF09JJxaMhhz5KtxE8tVf1rPTqC9sWpXQZ23AFubwc21B/dCu
8ErYleWbW1d2IeJc3ufwYadGNcTVRenRQ5eeCTkkXPJ34ktp8IY1dabuOXOLlD09
gDG0++HBqJf/RxkA5DbgIHRlVXH5ELHpnA/eeHIzoH5I9J03iObY2DZb0moPRWAs
BhfNI42L7X0JG6RS9fmYqGGhFT9OwqI+AnWfhGoNizqG6nKjUBPNWZjgol7ZkJ2A
vmz4XC8OM+Qs9ewSnVo2wRwE675OdrtpstDMswSUqqb2Op+QTgmsZEX7XiTDpnqF
VuZlH95zIE5X1sekcUPx56MYK27PRhtyjTmP89dO2fx1ZUOj7WVM8exj4eo4Ogyh
9SvsAppSBS/boDaZ3gWCc7nDVVUGm0BvlKyuYmU7tkQsZClNHcOYkGtKNoDFf6af
bDCziBC1vp7JDOhoTF2CarNLaciUxXDzJH+cl61B24ZVSzWcJEBvPf7wT/OkbbHC
WcWfYF4sLxULgoGyRrrZaWKSyz1OvlY0rtEqTVL+y1rpAw+uOh6bNGimUtVWtS3A
8i+JxC4VPaprnQ0uAxBYpWE1W3RdI4MG3XJkcbHBT/pDcjldFw09vkLTB52XhbLR
+CVgB7cQY1ABPCaHM0xj+ak4TEdDUA8Ya4wcWKOYWegkuhRBzCP8ZSMMUgC+47Br
4i/HjecJcAk1v8Ak+JOETqQkxggMPOROp5hA1sdbNJkhtvdbFjkX1gEpycBLf9q5
dxFIwY3gZtnpGPZDg94b/2aiBn5+7feV5D+hpUykTlwNTKD2eZU/adoLh9USiXv9
mw8QA0SbH34FzgcvLUs4qz/eHOnmGfy5OUe6Mhq5q4l9m1PN31EvzwajK4Sr5kqp
fYKNYIwGpwte60monMtpSuLpGPt4GRtDlgCPbDMWXHYAp66Pccwpazkyjl6BQTGD
qndPdjzt6YG8OrrLWf6Err9LsXAFKlNsmGgFU6LwHDiZ0t82RuX0Xu0uELhEMVD3
UHd+9ecRmLO2VlDCQT1ndKjt65sXYaoNXgPM4rbyCNWNlv2ZDGtvWS2lG0hhq+10
C4ejQEN3Aw79P9G6XYqxWBuBiNB+h+Kjyk0uQuPcYCqNjdLGYpjQQKJaC4RMUOO+
D8vBzLSlxO5PFmaMhG+IyFaKN0rdEXq0os+hr/M5iajVkTzDcuGGI1kx3TbxFNqL
xnd50E3eYYjVagkVTd2UIkUFHn+pZMdIiB11OAmUoM6rLnqQqIQ+i5KukzKsvlMJ
`pragma protect end_protected
