`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iGqvkluywTt+OqyBc8bttIJwpWwUd2qCD1+MxYPMFB5ZiG+b+ebE7lf9NUiUtUxt
/Ym1/seJ5LlODDtc4QLzydJNlplQE4/RpVin2ujRCnR10p//KeYddlwhvZPpwK+D
sxK3Hm8GuLoLWLhPq3g8eoo4MHBz4cUOv1OmmIbq7y2PN7zpVHrQokI6Kvg4494G
VdqYx1WFeb4nf4ylR6u6zg14H3vFnTNl3XLrUarR/P5aeq4wpmXTKzNmN/WUzdcT
nWLg713To0hIwX1eIh4HUOHYm3YIu3095U5Mp///hphBFnLqOe4+M0CPj0bK61XJ
wJIgFY8D1Xyhnn3SerRqcw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6032 )
`pragma protect data_block
9K9RBq177AyFqPfP1mjyAf6RmU7DzyYhiZ4k+hqcxezyM3EQLawD9PoB3wKFkrCc
ynaovMxUPjOxzsXtFfsC+mwCNT9aOynKNxbmL1auURIHmSI6qdXohFCZ3LPvL84i
iN3wc2XvvJeugaDwF4MaSKYW17AhMxmBH400LSSa6SrturTIasyhTFkgdAogvJAL
wvwO0XlLMB6vYDGzYPSFEWrwD1v0EsfvJ7vm+2yXrtTLMWSwe5e+oEdvx/DYy0T0
GPt4m80ShtM2E7DxhBiI+KtOIcHfJocrbrsKRLztuwTnJZv8dvHLHlUl6PBvoWOJ
0OXLGNXIhRZ2kzcwO0nlvsOQOxMJxq77Ywu1SbVJ4knvK/ElZxraQ97OGKqapz4t
Ypz5s6M5xLFnwkVYR9g/mUuAxrbfV9I6uQRboHjKZjnlzMupjlgPUzkg0rBB2Ev1
jIjQW22D1r1uYpT52EfcDu2CQmjFFbc4OTIRPG/jNgp4TKxe/EoytgzLpyrRAj5u
XfGn5BFlUU9tiwEIYdc0LGFB7PDtWJXqSxG18qtXwbVFkZgXNpUVD99eF0V7mV32
qKY4hFYqoQgh6nFQS8ggfuiEWrPHad9GqvbbRCiX4EQbc49zrH/KoVOIWTg888AA
qGetA1iuYfKdU/D41zd+trgKbdNm2F164vpRY9BD9yve7RJa6olnAp5DslZHsxy/
ULK5n03SC3XIkBeStA4E744bl7ARyLxbovjcEJuEtSCvPctjtQkwYnIWUMb5yHsY
pHpBHFS/v8d4MQu93oS+mz9OUnpU5hrkkUh0nVNOrAgID4kHKr7DhU02xA/apwtr
OcFcJxtryeDVupvo2gzjs51uO3k8SQmvgXgUxq4ZigI04EkUBAt9eMRk3Zy+Sj/l
zXkWoHJGRwXxK0NzfkB30cQQm1gWeYgXhqFfdTIT+nguNKS816I5bBbKgMDT84nc
TKYRvxdDunBENZUb1OkKyravcVVRAmZhuEXyCWqpLEcQ0rho9r+Oy3kogYxXD/mv
E3ElTcxyB2ZPbQ7+L7zMsFtWkc9ZZNfmSgsM20s4Dbo/8FNMZyjQMu4zc6amCn80
EEUdCkhhU/Pu6+KPjYDhjvES/8kRGTBB+vHT8u698A18XQlymAYUgWHlnUO3RZPt
C+8hQ8FVZH8yCXL4XZnPlzWnkc3hV8FGGh9nnkhgRq67sSFDdL5y5Cj6+3e61zON
c8WbioTw9b+kyS0ocx61urLsZxmcgHR+hE2IzQXto2hnBgkg2/SbK2tKi2dL8ERW
Iv1ddHKtZCOI6qWGvkOUwIF6vq2lHDkv2hGY6SdF2yODfz3hxxZ6l4z/PSFyTsSa
ebO7wb4uvh4++kfWYAL7llGgoSWEJQnDVYs8w9fACS5nslbEnwfMsm9j8CajvZH3
D7fY8NR+oRfqqptVg2xn+jjr3i5bUSXTGXgsxE+wIVUnKQx4FERHQeqLPEDH+b/c
Xld7kufM6nMoZEbM7VWOn3+9fdqKQeTq8x3zm0aMzuEAkBq/cBiKoqd1wx0Aimb+
QedTz9KqLI7VG5xTA4Lsk3B09/aW2eriYvb2L0svEU1yWUk9J7WnGDog7KW5WKUT
mpj9FBf+uRVv6Z4ujfeuUnFEiwyVQKCCQ/gtV/8ueEBEDWKKRayo4Y4kJ81K6TMf
T0nXuq/fNWvv6hSqG5VHwJHgnL/tu3cKS0SvV5GrRYzmQuRcw8AtVxtH+3NI5Yk8
RwMqNI6+nzODbArbJc2UK+w8B/r7YbANk8CMk0c9KS8yHg8xkOlef55hu2hL2bOA
T80C08Mpo+sIAHP79gesPbVfqDa2dNmR3W+1/MvZOdnjwxaDVm1iTAOHeQy8Qs5u
73eVyOUgrR6MgrAjycjPUCevnz5mbT/RRQApcnn97mM81c6PeK3jweeSS6tY8feU
mYUL5QGpn198cP8Zmx7zyqw3rnp3g7Ri7mTfsNWtJWiZLfzp85NLfJHi9aaX2g5Q
2qP4kLdwaoaJpagQ+hFBPPpEkwUteBKTwYgku9xTje2RbG+Y4u0OnjJZrDRpywj/
IKPGCxnMNfGl/WPKo5uIQLAHG27ndZu2zLYbYBgdrHZELMGKsSrshBV3NNoQm9iP
UxmhUZQ9uynIz8BrggpgLk3/pgGv5+he4CvAz1MgDIOAPr5CaHdEUPrBEkSvMPQO
/JQAxLUsWPt4cImyQNB4sYYZN7nqQ2R7zepuTLXtJ1eGSQq1n5LcZcK/otiDVWcy
Q+5QmeKR9Lk4gEgItBNb12ir9boB/P2mwzyWQCCNG17j7NBEwINWu0BRUtulK56a
xf/CYNT+E1lGBXhDAv1yUHb8c6fLBIJAlycwwuJTkCM6LFEPyg7yJWmtXjUDR7kA
i+xJrNwILF8VHksjynpjWemyLf1q6wFCvmJv1WskbkIIeZlgM8urdCTP6jcXgarB
MVaCx/9b4dfd+amxdeX4X2dxkOg/5lD3S4FeBPul1hrkETcnKDQDPXFeiUIl2Xfv
7Xi3EMyNBG97EGQTwbrVySokbe2URVv7SPcN2u6N7MYRiDnr/3p+xj5pw28VDn8v
IhXaRJWba1HD2EPcGmk2Ow4guW2q7u8u0A5+vr/qR1B8UBKiD92nDG8+FP3ZZsjf
XKtpV829ZGxigBr4uFZwhuLZG3VvHq2+YPnUqAbjgVg6LU4Cce5XkGA6zeuy6OlO
3z1FFxNwvmjunZDHW7WGXfirgdSTSpdzZxAQI0oHS05lwVCa3qRA2aMUgUBeUezx
IzkYCeFLKt5mZPUkGxqBbOVTei446YtIK1n/IgzdAZYLqoijbx7FU2h0+Llhe2AC
IdGokGcppW/ZVi1ku1wpXwryu6vJ6pEBwHgMfMuYetbgY9PqKyutWQGhSrwWzJzh
RIUSvum7XE1XztiH6BCPSAZqgeHRciBsF78j/8OFqVmwxtO54KvfBZknHRRnelbW
FQWoIZ/Qp5J4Ywph4ZVlxRwvWC4qy4D4YEUxCNZJGrEGiBx8waAU2hnFCKYIRkTv
1CUx50j2KKVWKrZY1oTb96S++aEuXLXA9Lz8kEZmCH8b2L6kmKXRDb2sYNEf6utk
9iR4JppFp5tq5OXq+K4A9paP/li7n65addzl48klt69TD36Tcf12tdT2kZnmm57/
tTpu53BqUle8HFaQkrs7WzqW9L96R0JaYMuC66zvL3y10rGJ6QJrk9ehMP/AEE1m
fvV0MPoKeC8nuNPqqb708DfpeN9/5DRrniVbH7czifmGAPvcp5rooNfTd0dO+aBX
iJyfTmvFdr9Dn/IdnY4aRR7CwstXZZt+p+Yp162naJDw22LMDpU1/9sX1bHMe4yL
nC+SwEMW9xNaxrrPGqPw1PMznzVbcmF68nuR4K6E/hBak9ufLCBijZgiBHbA9n2S
YoaNEA+eOPdP+UnbpdhtSUImZRJk0iTTQFMTF87Qnj3bYPLeGZQSk45o1va1M0l+
7QlGQ17yU9JGaO4sslVpPr8y3+tmUMag1vLzFHutl77cAcLg/dnrUqIDsnqj0BDr
S6FEvk8dVOTkPh7NEA/rnNdDiBpn5XJaghKNhpuaSJrI2Nl2jS630uCFbasYty+I
qPNYM6CbCI1U8mFcstexfH9L+vEiGy/AJnzO8vbjF+QTyqvA2TQD6OTjDOczH1W6
9ypQs6vJcZyavuTUwAlvgKMLriYl6KOTRftHZ7eMCNCJXEhNm0wdDS2KbDc2zw+s
pBrKAn46+phc9eDZqcJgJ8Dy51B+PA8o/R07Nj0M6ruPmRBX+Sj7UVZZelvMWVrQ
5F/gkTHKalq/z17/p0JaararSSW8dHBvaAXBF20Pebseac4GeP6nA7FYpNrMY57P
5kIFv6eSOqtfJgZvo3BofprEtVDRWJGHh2j2NSacrPorbJIhjCWbgMJrFzQg1t0a
eqMVjKtyejgaac/gf2z5B7zYfJWuVLds4vlEeuCbiWHNcn6sN4Y0sM5+aUe4g0sD
qy+YmhHjLxifCyTbDUl+C2ngchHqxQeb7CxyRGCHwpZ4LJ7ZREO1OZtOv+114bOp
7STrMKo4m7wKQOEJjIq0781A7BUCKDG6X0bxCmt8ypWm1K6ZJcrRGMZDxvP/KBRJ
TbYqM3jy/hkvwXlWIRqUfBAA58kv74Q4NM2OtZS2orL2lgz3xiX+lQmluwND5c6n
z3odkXesZ1XTsnOxGjDsWHHkzctzRw8c8cKbMis/4QEIYyrS2yhrIi+HihfWLjGQ
AtNs40CnVmD+i5dJAF8y0RtjnAo7LjLcpG0CJzXbSk5u6dCmOf3jC5DjYDcyDqcz
8JVvmHHz0ulcQu4gTVb1U29Vb1ODZPlTFfzJV4xYkVo2mA18xVO/H8hZXUfrfQDj
YdFAYdWV7uqfjDWX+7jDFNit+hsZ7Y0uMhzsRIjslihMfduuO1eKAxv+fgT/sIyU
dOoIw/4RBcc4ImjrcUw0QvPxLP0x1x1FMnhP7ZrLwOf2m+NyW/XA4au/7RP1UP9m
GMZzkCgWN38n0w9lC85OqmmopgAY/0Bq8UFZkPhw09YLYmqSJSIe7mebKIJtHfQ6
XiH7guf9oTZ5kpOqhdCzZjflssfXe4kVuMeXHTbVqKpZl/RvVvVBu7cai/yjhVq0
fHW0bx+BKGBgYYRKS3M0eykteRx8lf8y3CiSmEGgzkdbwWtMCltHRV1OUvi1ngx5
by/WzXrPAOwIR1kBRqjgNL7w9Q1G6utymjZLcdcEfvsNE37tDNfjmMLVkTK7ndRR
5+LCmGaj8axd5qVHYg0sFcgPL5Ig6BgCxdCuCrCSCyFyIXVC/FzgNTbmE4ONnWNG
2IdvbwZZvESC98EV0R3lfGJKrFdHzvn2hzgIzGmWYVTaxvuXJ0NIwiA6AZAZu16A
DqlLRDvCA9AO6UBRhns9lp7mLDtbtHBZkapFJ91/Gu2onDXKsIq44YFlCmhcrrPv
QHdhM3ZenvP7ZEP3olaS88m2NpTgm7ydS0KCFpUnrwHW/VlQ68IC7Cq+mUj3KxrN
uRtG5jEjDwNH8g9bfe9u2DTU372/CdghxZvleyhlIYL3UPlwrnQeo8nA+Y3Gf9/2
Axgis9dojgujcDrYZrD6sIBmrWnzN2CmwPxvhBDL3VwfQGFwdBa7CjuNnbKWqJqS
Es+MH+xr18GnQE3wQZkBKwM4jXAIB7y6afM0Qu5bAJwFYMV1uh2JfOSBnKDt2bgk
HAkvJVRNcftEoGM+FK1Crw7xzqAe5QEwJ3RUka43AgPdOST/Ot5yPsKQ9jE4Ak+A
MmoWS7TUCPjVxpjkhPGiq+4DD5Pojdgc/t9lG/8diBMLv7mGid96hrI4ZFQD3G2V
xH+QnKU0qFh5BCf8Ow4gFZ4uE+WfrPKSQxEghioDN4T37yl7MgcFIPANt3on40bc
bLXgZHH+8mWkN86Pouv1xcTN3l59cpE2ZtKN5Luiu3bsYWXnvYl3RbudkjBEh4bB
ALtOgn126SeCTZN+LVrPa4Pr0DevbbpQN955O3JgRPo/vnavlixmgR3LlT+yq8co
cH9OxWzOk+hFMlFBweU8iaw9FrBINgtCebp68mMEJWYBtlFhhG4QTPW3h7qjsLWB
LLeSnR5r2S2HlX6EYYiANwEgZnqmCLaTVa3IzQbUrUA//bqdUdIgHC1L4J/McKc+
64cCpj6LZobJvgNE92Gl5k0FHMP/umqy9QCloDTOueQeYUlhtpo8aLQqXOjVKaGb
mP4wyJEf5llVSYnPBlKmD/z3aSXQ4Ml6ZX+18j0GGi4ATJKA2RwMr2tVY2cxHQkd
Pmcllaq0EslzOHZOUTYzvQEzcszpDC6smXeI7Zrk1kYCelbhqz5uLl7p8In3nuHY
1g9coibFhz4T9UU/XQyTKsv/5lCupg9oeAmISLsn8GlhR9Z+EJzC0mZ58BmOCDF2
5AToK/C0BM5yMLNuZh5Y6QRfmhfzgT3vDuLR8EJti0io6y2VwjJG8w8Ny8IaeFco
EeZTGkyOzjc02LMFVFM2J9ux7keWg6hDcBS3bmPRyRgamAH07dx9hTxroZseYqKh
y62z534Y9IYkHYgkRgyc2wAws+dhnJRDrVnYIOxmgvOHGbsdAjcpi+wr3soWi/P/
X5fwo3O6E1/5ySPidWeFtm3mmJFz3Ge35b2Ry+vEvGKlZ/n8fafNnZt1Dllzjt0f
QvdPK69JicJGhdhMyrzu2G+P9v0uS2z2i3ayIoUSfMH8oje+myE47dAsyB6CIyVe
sNgl/ICwVtPsj09BX5jqeavZKVeE0CBb4oolDH01pYnytq/7/y2E8rWUswrXojk1
S7yuS/Xoh9guvWZgzKWyt0vsLlI9SB+ZEu50R3TBa0vbiPGMkepalPfKJIzV2Xj7
ZxyfZrwjH1a/FswRHJZdUxy+kKJYgIkVa23xNjH4RT5NDQ5Zxptug0a0xwseDwS7
VHdaxmXr8pxSjRBTyi56UYT2v4FRgSibw8n9m1U9uO3qxsg+nB1qFMMUE9hkRSQW
N9yHN5NezfaKAPe25Y9hChPFn6OiocPWj83zd1Znfojg103vLf/VR2HxA2H2hwiJ
sY+IcWpd2WRYzsqnU+WOutmGWgLy2brJOLwJWxTNurqIIARmLbCcVRse9o35yuQB
+FwlKQ28rtvNSDV38+DLdJ9BKfgcrswKBcpq/7D4aN40XTbqKOU6C5sbrJvCG1X0
7uOIpxnzT9YC/3dH0Gg00H1HjeZBU9eGmCluEyTUnoVwThKbLZHnyyX4e8qyuiVs
K6sBRD9o24tHBYHpZzrpkEldK7XU5K4wBERLr/hPBDbqbkGaBmF/vkMf1D71S7wA
9PYx2fHCrE5nAyirfz1ZUIRzDwFsKS5MXAMPW5bimQCXy2KMlOv/CcVTCvN/3zqd
6WtnjcrbBF8jyRs0t0OCqgN6gY/gJoA1KdJqInbokRW32Nrv7TcY9xhFL1CKGoCA
Gm694BAEN4OaSYurMsfRKjI6bk3jDllcX5kZlH89eo8/qZ6jsWOKnqHpaHtv3w1p
/i+4UIRv3CAKqdbC0MVyHbcarFlZx5ewO6nPco3lX/GJMT9xfOwn5Tnue0WDi4TZ
EvIfkbKPz08akPaiiKAO+bCKHk4T8+euroM0IaLGlyxPsDyp758B6oPRVSbWVI7M
3RGfr8MOpo4JrOPSSz5uHmxIWsFvjnVlk79oXClaCDIpvRtMqM2CVibHMlIIFWJR
ELHsCJydSn6CLpZFLo24m0CIXLUDO3PSYETbH57s4z/bkj2T/HnmTin9X4CVSK3V
eB6mJ3OZXMZyGXRbwXIYXvaowrZVbqEeweNYNx0Iv8r+1cj85icmm6lFq56lPGHq
C6YB/3eOYeyAxS5x1GnJRVu+eRdhP+aMiphstP8kYxuRAD1CxhLii0NEr5vqH7fd
m+DxlmCJwjOmH3+gAiP5vFhAG7KwjCaCWMsBcQrca2z+zzDYCx4afjK/vF0jCWHM
RUGLaQ4rzgnNTIvqBx0hk/kukHWMd4eUbZTuXxCl9Rwl9JY41X/nzhFWLE8WtBEb
aLnjP3l0uGEgs678qtgz+6KC0KOiq7xJ4QUIHqheGrsnHn+yMfSuDJIIgE1c202x
M/8NAytUjBhTv4sjSagoei4wCknEuY3YLol7kTKBqS7vVNomAy2IQsigA6JzIwMi
5EeXh+GrL+sW1czE60pX+OcJjwIInn8VsAqbkOb8w6v22EFk9P3xlzJznEsJLEp4
4qhWxFiWEAR7PP4bpCBUhsqZ8o7Wle1qcRGkAlOBVEFFeILzBt8uRWcViQpWRqGV
vQglgPNCyCnPUWUPmwdDIDhNlt+dYYQmyolaq09IXtH+pcd8J+QsGjtkKBbVTnsy
ngN+mEYiJ19dvcSt8QMGOPYviN2O2ONFN5L6inWiRYff7IA/cF1xR7AmYYlUyY0Y
3kAt/DOYVLHsXUpup0vLx369nmW+OI/4QABQt9H7sAbDwBPgekgE23zZvO8awIeL
Y0Z4KPQGCk6VAI6UOq7Ql5jNcPdfiGElgOuKDpsw8LeaZhta0GgZZVwvF/Zlmc5F
msCg/CUxZSlF1Wi80GPBozHvDGO0W9GbQBYM8cro8Zk=
`pragma protect end_protected
