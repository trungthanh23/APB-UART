`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
THMXMdj8EBXXMSlj/dobFcLyestMVgGSafjxzidTiVS8K8YWm/POJScR3CmGMOcB
M5yWTQyiST19FiNsX/bEOP7a6QDhCAUtI0HXiZnDB0fqkCk9ZI84dy+6KB0ngjee
KoXrwcalufdHY6pxYHvIh+ExYX9R5ziys9dK77h+mOhW/tOEugfQiE3qPmCtc0TJ
fu4GLPmKEfgXh+RXn3tlxtskb0GEl87kNtstOgP9OyyVpqdBKpQhGRDtYWrUVY8C
KFOaCIWGH3n6XgqRJ/5HQPqVT108UwlHeHRa/TRv9n/oiakzR2vUmpMjXkj654w0
tSa3HgT15Ggo9J5NHPw9Zw==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3360 )
`pragma protect data_block
sVXD5gKvO21UViE7vjcVmefriKVEGLSHTCaNZo3FF6QLdYhGOCXph74xdCffhUSv
YJ0TIgHgAmeUyBX+WUCptDBozexC/sPTecvTaTbh1Pyd48FMpAgPDeJu3iVXf9Qe
Toxp9Y9kTmRTk9ayXpOQ3CH0vCfvtMGIfK/Mept4ILNOIyFlTjBgwQxndNgzfGlX
lWZLO6v8K8SoF4ivgPVjwmO1GR+LWJOiw8u+YUNErnf4io9ZRS+KdT+79NwYbHLq
d6tNNelT8s4ZfVz3PjybKQZW4edS77HonX5Slq9ihl4b+7Q2yVKyUASINT6aycqH
KG+BwJrkiT+fEQbcXsAl8TOrCP8P8n9bG/z/OhQkd86s1DGCCj4Ks4IK58bzZLqn
wWtHrAeesY1Xda0HwAwSkMgQz4tLKKYLWcUl1oZ12PZymXVnV1HsyZZfzA1Vz62i
e/tHeEQhtBY3BOpKXwBjQEsTBnthp1z+FkoNMv9QihMI/4w8lFyHyoJV4Pvmkq5r
JvlkoL0eggEDeJZRLA0fEETaFikPTsg/5+StQGvf0SIXhQAvqf2Ja/r3SaKfDi44
zgNSEqEw9y0dUm5gmkMgZCiupZqjpPTBVgmkKXoBj1u/MQv9gH6ZTxSDZAW2dtzY
RJsarxSOiHywhnYl6RlLpge5gznZa0mP6tBXMJLhRIdsmEoLgPrXVk2NkT+VyQGW
49uZ+31HS2MxAUkRFXlmox7rHBO/7C3U+Rz6OshJaPNpxNO0NJbTHkbcVPz8kQV+
MfcR2fvDuOo3iNRggngn8pI70ccUw4pgMVOsrB7/GDbzNewr/+e323aikGyamwCv
CGmi+0dubUe0D+NeDDrWsDAsuIZWkoN7hSTI8QU4jyh/HjESaFagYndaIRyINVE8
iHB8n+rDB3zodJhN5dl9EJw7HeLONkTQQLB42RbKx+wgm3oR8lQzIZy8R8139CWK
lvRZEpwWvvoV7shq3J/qvRMFVZZIHbNhWyW0/84C2MtwTPw3O2uCEWoHhFHcRmKh
MWcHnPd1zSiVAeWo98F3M2rJJNb3AO1s37fOcvpxUqc6Wt245xaWF49fAK/Hw3rt
fCnddFvvhMVApkrmfDwP9UDWA0YAtlKZUftExKDvGoPgTrT3NjdtaHl2tYCIZd+R
SW2iRge3WR7vV9gcrOxXXahO958Ob8r7oPvmkSHp29dWk4P+39HWyySEwQ3u1bAW
DkRpyyD+ObDPsoYNTld5Kj+IdBJoCS4pkyVqweG9JGf0S6ZtsgpDSkalDj3ucnvI
ALU80i6RGkmRKTx6qoa1bcRbPTl237Zl3GGEKXEl/BPkGq2Slt/kaIyl5GpZI9G5
ZpqA+n3ZCELXWh9FO6exTfCrHwbEKIJPJVWiy8Br852pyENoqmPrOa9k+Mu3EpdV
CPskI80qDq9aUXwh7jbd4lB/pLU5+O3oN0EEaBr4eOQ+O1WbrDiCFj4w54SyyC4J
UI9AKBMiK9/1uRTaZ7YFCKy9FVIyqu9tU6T4pa9rMLYW5yFvxI8Sj2woRuTUz2K9
wvpzR8JxhYvAxg7AhoObjYsUywaA2Ay9V6iIYuYpR0o14tXqzbjKdkGmTtOFb+i2
+zXraAyWE1xFc7Ov7Px9sdhKBdhNQlN9BU3thJXzx4/3j1A4YrJZjAeSlaaegCd2
u34Iv72TZI1XRupbkD/C4tZ4wlSXEWUesD7Wk7dPBePdcvwI3jfcvGHT4YJ2I/Fa
EvZo2yn/iKJQP6WBYRrKvZgKpVm/Nu20pZanDZG5QEZeGbcum4WXyYsNOwOrO/ia
ceYVDIJQQVubTxI30QDN9RR5VqZDUVAJsUQwAzEB5t1AaCYbFU+r1mezJUEMlCn8
nfce8wLKQlsU6sdaVIdNqGWlEejXg62OjN+40kP+sksgHlaWXk0L4z7hU4OPua2V
j1qC+eidMa6l4ry0XQgHy8AtzwexsPd/wvpJ9zqH8irED7klVDsKQZorDYnTpeGh
iCUc7xbQJmYnXvUHMOyUF+afJXzMyFJbz/P8bT50fmsgH4Ohfdse1oeUdImSF/Gu
7cp/Wuf37zJD2KSfaNBmgQJroFJz7KG47om+xO6DgZtsDlbD1ue8Hta6nXcsx+Ha
fhpfZrLuIEi9HxmqiIEo//sRmPDb8d28Y3PGsKgDcjovq5xxngdwEjjPLCQYy0Za
/R8s5VoyvhVGw477Fyl4gsEvamCqyrCU4s9AVysHdSiFpFOPS45+vu4IXMDxixJs
pHzpMofUNtmieKjPxB5yprilX5KcqlpMp9lkTJnxX9vdFV5kkGXTsDhCwY50FvU6
wXCXqxjv0ADXq459YrvMCBp2ekppmbPon5CesYfqb9x0593U0yKvoZfDqWt4HU4R
LoGNP27U5oD4LpPmvIG9RhqkpA/HeVvMHyXamgRToPITGmfgG2Fmn9u0SJvZQk6F
zCbn0dV3kncOl2+wVRR43lSEl8rnosMdsyV63DUf2sUeBkSw95QyGCIXgggkqf0w
bEF1Kmrm+5aCnEWlE4oeJHckr4kPOIIJZipooNHVGFc2Jl47lrS3IMlEJAcDS32a
9RAT7EhDMrhaXiUwtFemLayo3x45uhJVI7DZaju/mpcmM2C17OLJKyFolLviiLm0
QwqNnucdlvKyEuCjBCFzNClQRiKzZPNEQwM0hTEtI++m/g83HarTlre4d4YY2BwG
e62P1TN7zNouahWHA+4V8aTkzjJgFI5Hp0o3XKANJAWhbXgh4tijy/VtGJSE8M6N
870T+2BM6cTMDolIheKNya1IRkkTWAvxyITQUqb2WnQcRF6CusnVMxLtv1UJDUrM
3xau3TLITjeIDSzkmpNqH/3MVxVLaE2p5MUAg5xVhKv97WdtVr53njiH7qc1OmOl
eH4JWd5xXiy58OZ+SzXFT1JA5iTulnQOKGRUSJUBVz9lASmZN4Vzm6rE4ctSmJ73
YeQUad4YwxsKoNpE41R++epPjFH2rhHBOIWE09/BfBi0lLhDGbgpMHvvaGwqYTeJ
Ib8X2d1YqdytfLy0Bpz2cE+UkcPoJeiffneNo9uPy65Kh/SbKGUIVSYTCZUW5Ap1
9dz5P54z1L1XDXVi8d/uU/7NaM1HXoIqJQIwOTyF30C+c+ENQOVtBfrddEnOSrYM
brEilz9MLF5RtSHuGx/MEmclWCdDQ0+eUXLXtmnm1XF2OqdWKw47ZvAWJkDaOSya
yRHCAI3E+/yLa2uIwuMHO2aEOvixzfkZkKtO9EhN/RiMRC1hYGb02ZB7L3IW8EI1
yw23bSu8lNazWQCytvkyBSvARIdrjsnVkiBT8bhdQFY1UdWr4f/hojoETHl9g/3j
vmOt2K586aAU0HPkQiqX7rkvJS71IfMJ9p0dBE5dh+X4BWmaFHol/NWTZoxHZwz4
yrElj/6ivAFcei222d1bk+4CUcxpB2gujV8h6baoXQzHYj5v3/lBWRRKj4QL/Le0
b4cA8WGWOixATEIfztUy55+STJxAND7SKTLAd9nTNoqOeTidVhP0MY9c22L/TSaP
47ELNzLlxSy4z9U1feYcDm9EJ/2g8/m8OWoAALMM2MbvgO8s3WQI9lVJW3Qao78U
UBPH9BhZw/Windi3COL5QGMORTIDXWirL/iAWoPIqi6Lj/PmxrbmLfdVB246ii1+
jOq5Wq7926MTgGC9jv8xsAQOPmv8bAfsgX70ll/iLzA7y8d6ue/YM/SHe8/DC57m
dkYN3J/c/KV5FZyvPOnjB/wlnXd8/biBqhsVBIbUjPzAy/IIrREtHaFnLbyK1m3z
lb3L4rUXLo1QvQxqHysfvA9eCW4p7APTQvHX/hILxjnUvOTSnpSUuH75Vj8gLtKI
999woee1fd742a92d1+1JWJhb1dcJBdBqXecnQBcUDJRODi15o48pF58Q8beJyDP
pmcT7hEpX7jl35Q+1kndJ20sHF57TQLb1RD7KpYF4mGdcHHXzBaflu7GzPIlp781
NIauwBwHy8ruysp5MV1IUdURt529qxRAA5aSysfIsDaJ8VDkBLkcF91SpFF0q4ae
jKUZJqmkVuOFb03D5jJqhmHF8Hw3i081thsvFeSv63YeQqRi4SoPv2vMDGwszX+m
L3cw74xhNGG5QTni0mOWMtdMhjWXI556YMnK7YT+crCObjakMhaNhjjWcgOnr7Ok
zO/rvUrQLoMgkNip34E/wP8RdqeHtUyYM6/8wSMmCCKxh1qnfbsnyYb+cwRZzyrE
34xc25lszynUX1ED1oUyafMdYTZ43ZnC+EVZ+E2T4ttK6/LVaLpRnDFKx0Lkfhia
o0oPpSKqAwN+sDUl46ILVqeanDpLifMhhLq5kbdR+QFMHCeGYoL55F9xHjHFZHuy
SlSmlegbgMohprB58gyWoZ66lJ7xEU15Ezf68bRVVZpFAkTfPv/TSiRp2i94ycx5
M455QXXsS889jTagU0DXKJ1a9TBCAuhqfTB0guRb9sIUW06C65YmX7JBH5FCL68+
`pragma protect end_protected
