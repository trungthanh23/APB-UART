`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "10.7d_1"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
h9kr7Tl/HRJlhIK04LnJBiGCNDe3zxtuPIoqOHiZZ451Ny2rAWMRZHvqMHN4rpqR
X37FEqXrwCToF29jrEHw5IeeYNEKbyCImJm41bMZdfpD/FMjqoFaDKUJmp1ixCYv
k0zW38crmFxo3gEgTT3vSLYZeTv7RBoH+XplQS9u+BTpCpHWd7cXfnmcxXXde9nZ
3EPs9w+6Mjx77qmeymsDRx3vmmSuA4ZyfMxDNnx3zoML0wW0ayNheV5VRa9HZ5tj
hgcD8HWGy2zOtbsIqS0da21KC/ksGkwDkKudgJTOX2NmnECWl4pWpIupWEEsV30K
rw6k/rurfl+dfH7R82Hz+g==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5520 )
`pragma protect data_block
TBeC1fAWzGC2YFfxHi7/662JfttX+aEBavaNR8s/oVRhzZTS7Z1oNZ5TEgWHWflV
6pXVhBGbc/P91OsRhyOgRq57U0undoA5iBweJJeIU7qqygv9m6I3asm4Yigy3Dwc
2+DGSi8Yf2Nuf74d67LYBV5uFsUEoSHu5IAK6TRohCTX3vacfiaZfeR4Rj0o+bpA
koI07myYrc2cbe03u70EsJwSK1G5HMl8mkRl3M278+3LXdHSxaKicKfnKho9fMed
oLuXTaPYxGAahC75wXWFVJ3HtW6+LbmlKBRuNh49ThjZQpAn0vV+vA0DRegm08+V
Xw/Xx4qDa70GjswddvDN7ZsqTRL+PcAfgAIvmuYkz/ywOz0AFOGtA+2pV/LUp64E
kwQnOtw6hWOaFCudtLxyDkxSeQkIAiS9thfutvbMeJJ1oqoWupIjUNsbGw7H1WS1
mhmbAJJq+bIbk/wW8eSk8xW1+/kIDi8MGqbguAzYvjLZBRLJX+aPilqWWnkAsaHq
zRm3OAcVfM0ju3gdwowBb1w8RxWkU+N6nOyLefr1AqH7GYqcy1e3CJ8bObHe+jgT
rJCSQWzpsZGILT0vfSBz3pJ6q8Zb23AhTYVuS5w6tZJE+V6sZzSYvkSCz7yB4eJM
dCfpllZDNjvNzOJQhPydVLG9cVspOaMwqniLrLtKPI5TpueLsgP7t5PeajDkNuhv
szVx08cycopE+LIEDmEd7vD4O7sWGxtfF6H4t7WtyNV61TYnlIuANsxz4qtER/At
9Za9KoA+TpQtdjMRpoSYLkVdyICrFoakf2zQA4UADAwcmMipK4/y5YWbk3n+y5A0
CirkTjLDoGeVbUlIQ6RUzd7qgbNZdoPxd/2BdLno0238Ot02LsmUqksHBUmbl3Hl
An8+MWMKlTML99G6gZqfT5rH5i90GjOEDL6uEOWtG5riyOxsxHVzEUlpNpeV169b
P4CyarZhe5RP/VttjMWUXu/cyyEft3+/UfeDd2Ded+qBJBc7kIBYuNoAMgC1l1A3
tfgeU66PbV8FDhW3oigEpzq1KrpkC5l3ShsKO+0VUW8cl8e9apYbxlBFBXDBz4/6
EXtuiwN1IGdbnSU5eSCsv+22BS6AcfAPCjlqm5PgVw38CIlr5Xz6kMIoRtFAFFBm
H5V7xnE4/1o4aeWk83DYZPTQdyXNvnyaRy9McR7foPm6vLdrH3VS91btCRzMvLD8
f83xJAkBO1GXTNQctw3vtAbaYZUj/KRUQKasCkqCTXij3N7BV2gCc7lqSt7HsZH7
o/+9ZX7RmIak76KMHQ5extlTWQfa/rXzf6Hr+xC4J7wwPS5rAFXklRs6BSUPJFeP
LCZxyQE3SQH6ce9jJXV8qsJsXsmv4eSm4+B7ynPcOk8Gdv9HzFnRl3qI9UpmZJYc
klO5kAVoFB6Pa8Ku/tAxDJFvB1zn9jJButkA7kNOfWjhi68WPVfna//KofXpQ7a6
gdssEmvCFokKgAOvPscZRsEuF8vTv96iIac0rUz7sUcqQBDf551iaYXY+7Lt+OKd
WstsEHyrfbQNw/fhMdY5Ih70w5oPfMkTLpyPj5pZ5z/HGwyT2Dt59HeZNDNrkFsm
pQiKz+y6uefkaHIWmrq8K8LIZTcjBtWAKoj4NOjA/8W6DcXTAW0AP8AgGkflQI6a
gRlVzff31L4Ysx3Mhw0HGR1SHCqTje+Xj5rLTI7SLIv9lXB2dL+uuiwvXXYpSI8b
3QQaE7F0U42/O+zB2qc1no8gdeCITQxmWCHsx3GonO1VRzX/FtxqLQcjgAew0GSe
1IQX9Y0b56KKZnYm3UprTWN2OTa1IY5d8wo0868IDKGok2WMg/vqkLlBCID27tDs
LJFqLID3mTtiElbUXimu7C5D/qPMzwFA3mrmlYckBtxuGqmIFD9BZXzVSUjpk3/B
P0UgLbKiCljcFrrMHi5oTsnQGaOmaLawklh0tItfwNskFqktHesUWgBxFdIRazo+
tz1xeAMXUcpMURVHgW5IaPU2aItjiQ6C3gLx7fAVIhWjz94c/sylE0rZoTosdg+G
aImR16N4E60zo9Qn2Zb3YyjSWQDkWbBKZeDIN9t809Jm27K4wbYGTDtMiSd7Pf6v
L+7A02gF2ahLQmB5q2pPFs48s9o97eeqZff4wFuisehSi8dXOqslTnHt9Yd/C4jL
IVKjIKDeJet6R2qUQWSOxrhrPhLczEH9ClkknOzM/C/eCRZB/Ur0O9KdoD3wJrTV
msazk4q8xkLHGrwbRCu2x2fvnImhb3zxiPt9jHIc68y2wkVuqtH7/RjfkJkiJC/i
4POqYb77zfXTGdMulEx/Ku6vWbPRW7hFo4kGpLUE6LjiUkEKPyC1sz0PVPpRbk+k
6cauSV1D/Bo1putHWSZfXfOviBd4ctcALEVLigqzl83mP+MljliIBIDw5/AeVKxx
hMFSL1jnau3zSEKx9+6Vkfok5fBnQdOAiMWA4qO3wyAccQZrRoU52WzhnzEcgqN6
0Qh9Q1x+uN/dLe1j8ChmaObB6QjLeRkiLvmA14tUsnUUAMJpgK9Tqtz1YHq92buY
DThQ7ON8p1Wh1etViX+LY5ycG66Zz3XSL71Vg7qGS1EdJK7Nw4XpZFcQ814N8Zcv
NSYhtU0HfzF35svmRTMO6Jhzjph5WEphtrJRhMyszoDj3jUXsKLhlt2wuj8tnqhz
l08dl1/eVCHfWqJStlUP8CZpjs9QRihOvah8tEFo/bGng399mjpQbrodsVvqiLi1
cECGZ+ZJWjRVJQgU+IsfYMLY8BbiTR58l0QICpF708cW78orc2gcHrLUcB+fWpyb
GESnrx4MSI1h+pSpiQu813HcrHQl/dVvtPA480k3RHOVeCFQlUtRTEj/2aJmJV9F
VrTw28utM4hQThwrSMIcFVry0KnJGUjmC+QH2I4KFy4bf+9Jjf/k9WOyU+7b4SHs
sodv4KkaITkG8LeBwmwxgEyM5KoM3mHdasUxAOzZcxirchS7+M3ExjBZMKZy3O3h
fP2taacxYdvMbrQykfbEeNwWbDYB7rGFdXMoNVEgsYg0JCCxilwkLdYq0pYhuFqt
VgBZGRe2zRITT7hzCJnY1dJJCsQYbh6r198eFTYy5U5m/uWg1WIjvH2vEK8KLowK
/lL4QCO8YPYOJgRPuOXvrOwmm+pgRGb7h14WBORb5Sb9PADBsLmoanMtGGjyhqC5
Lg6okCUJSqMB3aNke53kVXdbxhrs2XP48cDyxTAtkOrYXblo7Lbh3G54rcQXQXvI
VDyHRZRpi4zK/Ypy3tXa9hm02WOEwaF+jG9Sl3+iPjVQ0EYXZq8YTa36MjZTYdR/
lZ/0RzlSUHupXBk8UBAhVCYk/gMqrD8FND9mHMpkW2T95XzEFKpLTyZtPZ4PK0Un
bMemAzofq9vz8VxFTe83YHqgPdpRcoD8KfbQ446oRlr4phJRu3A1yLHsOwjR6nHm
jITjjD9Odvhnxo55qFvB0cVTl2JAF6XrBX5GbOb0zelROvg2GXx8xPhsVRFrkP0Q
m2sEDJK5urFsS261Xdm1BpZB3Khoheg6HAw3IS8KIIZDIlPXHhkO39k0rDIUh6dk
yP/aRZ4i3SbaSTjkNpuWVnbO5xfBo6Ru1ul2GUSu+utXnHY95Vaa9lLqKi3CR9xu
OZdwIvw7NTJKAuRMywsxrc1wpm25/XXjru8ni3tHgSRo5wdJYbZ+vwS4vknryULP
2JnKGpMQuo6fUBqk4nIxnYAulioMGMmrdJEXTBOTnZ+ljyyFjC9dRZzh5+EHmk8U
X4QhJ/QiZeFyjYrmIGk+IQ5QdDB2QkSveitMKi0fkhhtl2YxrLqZpDoIy1rpwepk
3uVvVYuHxKjlgZocP6RCe0cHGtoP0ZCFj7+4qNCBMBhxTV9Iz3CglvdlCy7YHBKE
SCGPLb4LIikQba2AdK54YMxQV0Pb+1EUY8vwWEYyTYW1xIGc/5QodMJMbyOVzWpL
dD8W9mKalXr9z/Xs8QESbh9I675cA/atZMZQN4T1W5tyBVgqb41K6X+Dob+f+U2H
UCXOX6QTTDBQXAYErx8o5ldN5zkhFDarALb97lrRPHUFR9RPZV9+vNi1oWqN216N
vlO56uOdmCUOhTLkBwvQSR6/4NaHjqFkvoJumGxKYzvnf+30i7x8cUV7zdZg5DBg
i8+Ds9w7hui6/HJTNwfiIFZQ4lXcHgURIhIO32PbMnvg6tYK1+ASa2lLlpCHLVH9
hbJ4TdkfjkRHQ96E0YozRsSzgBaVi/UeWlBr3hoO5pT/Xdv9zbw0wypHIKdQeJy6
ANIbF+f23MytmxHj/qJtc3srRRvLjMNox3VhfUrseWwYvu58YoyOkuqMJ7hkoupz
zzMi2W1ylna6vvHGwGv5AXHWi3jbIkhzIfqeGBlTOWuXZ9sRig5OPwAJS1NlmchE
MLxtroHhF9wb84QB4lkX9uDfs4Jbuaem52rNDo0jmPhjtBcIKLNs6QcW+UyQZOkl
MnJKGoPZZiCW4SyoJrkqbdVYh9SsHv+kCVuWOYXjXJI+IarBsffva1/eBB1QqXmY
NN792gH/nWUGsAvCVTSAkg8Bh01QMp82gszgGAK1YrRVAIajeHh8csKtkWleQG8t
rvsSe8qcMmAR1t6/aZNNysIDb8XlZj+ncFUlBhFWLZUcS0XSErF4mx7upg+jLEWj
g+sZr4i0PcTjdnZ/ZE+wERSwf88Og+Dedip7CGU7koLHXQ+nN6ltifD1dZdnma6d
EV1Hv/5yOEdwDqWzve41WK2kBKpULdY76lXZVEPrgL9f0yl6yCoG20r033+rPBEf
IN/mQ2MwHvI23+tPKkLAiVWW9LKlYq1BPybfEfxGQK+JfZ7ny2aLzgslKHQz8T4p
d6l0PDlQ+Tx3DFDj43EBSFa4ODzmsNBfDw8I0LsqBluKHDZMwGQGwLBGMY6VwJCM
mPo65yUior6LD56JMQO1AKjhBYh0PGn9kxPGcpw/iV7soFWp8F3NNp8WtrCEgcBl
fzTpAkP0WbrwrlzoAJ0ic+6J3b2VQ/PPUwCW/fOUuZW12TmA7O+XP3LaXO429QXl
CS3UxjLCWb+fwH15UeFSpg0q+BvassVGFoFY8TtMLzXuRnymhYyg0EGcZ9DjKIEd
SVMf0CMpMMTbZFp6Rl6ZVxbEvSw6vqv7e6ic+51aMzJSIjhz1odcoCkTSVLtJOmL
OTJpBm1pL2OgJt/VW8raKD6+xLpb6cwL5USSyqXAEd1Eg5D1mv97nC7i2Wc+6DX0
usCaYwZr/rYfkGpb1TzLokBzQpbJbSEH+gUD/banwlb+FhhivyZa4P37HnlM7vad
idhfQ+mBS42hhLfWDhV2dHUgXFi4iwboXQsWfDpCbZLVWBXDo5dMhXDZ0nBeOrHb
q3XVbcUHyruDsZMT4wWiKNLnlH3p6Ez8kffUELQ1cLy6nrvVMAMQs7FP2i0qNJl+
EwA0t3Yh1f6NdLyj0lqiScGbPmTfnjZAtn9CkB7F99Qt4/iYwMxyVUc94Gyu+Hx8
8yRnoW6a8lVp4GS2PRXw2XyYBbrQDslkBJcFG17Zw2OWzBtbXP9/tKIlCRimP4hh
UD7PboH3Po01ODCARp1xJt5xpPlPExyO0u/qI3VrPZQaHGuJ2Jg+F3/uIK0yR5V/
mD9FCCcItTVK9prWZlOLj77gDSCwmD/DfBBwBWTxzSaZBX0C3NcmU1zVHR91V6cD
deFuhXUCFxKJbDuP9LXCII89eV1Nb28tqdUDX+/U0QsmuidyFWblcuUXX79eVL29
0IwIbYrsN9VbjMm2eRxg6gX8ICe3T1HFVKThEXyGnzNDCHA83uE6Zet+D1XYETTO
1lD3vPUHKXKSPKl+cvAckae6Ts3+7KXF4zJzD1NOgK5NUzm5M4u/H1rBNVYaYyKs
4iw/HqAOJYfO2uSuUBGa/44qKYKM3TH8NPAMZNNiYE8P8nFAfAISbXYrzdZY0yDM
cMYpvgOVg9EFIS3NgJmamfC/uaWWqE015RZXByFfUTWwhoFxXXH0d6whSoMnanSp
2S0uatuLxgNVFqru148Onc1TKDIoDPEWTbLO/XvR5UVH/xO0kxZRiEFOeJ4lg38X
rFyZalC+vcFcq13NgOHTZjqAjzMgtbgPssNRmLAISKxJXlbMWeXZllgHITh+y9b8
jEgOXMufeJAxSCOj7KVjW7LOcxAPfiUiaWnivknssvZapd++lM2G2H/RvjQYf42G
c3BTI7sYT6GV80pI1RRM6yDzVCtxPyPPU3L8ygAJGEicWnx+ggIX5MvoyERhcq9X
d1ZjM5Cbmr9CR6+U4cgKn7f18Vm+tQ12D7wgRED/NI5b7KDj+I7zW5jwnXjfY1v9
nXZLgI7udmQkbqXQicenBXCIslYl2u8HMYZIYE0Zy/qh6QT7JH5lkHRUlRa0Fm/x
4SAJzA8uQQm+ErpyP3YH4xt5s6N1I7tyJ1O+RXj8D9G7G3xXrYPLpKcv/hRGDdYO
mE1udLEyhYNgMc0npVWA/lJWMpJqzJEwenC5c+l8oJPlt0cJ+8lH9uUxZignP/bo
yLWzHCMZHcTiwMx51n9S/WuQnZsQ2IGtAairQotKMNxvex9DaCYcwq+aZxja4VyF
mm58rSN5BhsJu+lN2MKZ5pgjk2QxN61vKFjc6k6n6cRL7o2tjrJD9FVw/uaQhR4l
/QwDB13pwmM7LerGudOg1wQIjEpxmgyOUPereV7R3m7hK4tN5ZjrG6AldB+JzxdX
0jD5b9ffvBk5xcOHHP8DjR8fO+LRxpNFw/cikWgrfI6JiqIyhVI6lft+IDHXa8o0
woAu1JbjO7hx0yMeDWDUlhrzdA0LWtYtCpC2exBjLrmmbDXbNfTo3qAojeK7Wir5
BbtJxOWU0fERxhpoMTLzBoqCfTmz+7AVbQHHWaqBXhxoQWcuKppkF8he/IparOop
U3kQbIGBvCqmw4EfdDFmAYqOmifaz/F/iB4ZEMLHgUEJBw8NS+nE6cp+skeVruR9
zzQ+ly77gqpT0LTO+CxsEiFIuJMEqpVfJX+OzKx0YzDa16+svCAVYHCLVgvrQTZw
TLSGHxIv7HfSoigLSs0ufE8Ir4SD2TzmJScV3jS/nYee52kxZb7teIi2x83pA7+5
8ByST/BfPGt6LGxxS34I4HCuZhNcTEppECtt1Do4VniZv9Y6S515lTO5itryImt/
0/5O4QGEO4AWeVMVES80jIahub+x4BEN8QJwNWcQ3YBHW19PY2cI8/rEOpVx/Se4
XDkHuIAH3Hf0wgdUDaB9qzGTc9VybkMUg2nyEFG2gdH+8AE2OC3r+XNBxmVME29l
PkCoMc7mvJ8+7FptFrcdOKenlV6oHfOQiR4qwO9KxX61vb1w/xmu9kcLot7pFrio
`pragma protect end_protected
